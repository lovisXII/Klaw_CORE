module core (adr_v_o,
    clk,
    is_store_o,
    reset_n,
    access_size_o,
    adr_o,
    icache_adr_o,
    icache_instr_i,
    load_data_i,
    reset_adr_i,
    store_data_o);
 output adr_v_o;
 input clk;
 output is_store_o;
 input reset_n;
 output [2:0] access_size_o;
 output [31:0] adr_o;
 output [31:0] icache_adr_o;
 input [31:0] icache_instr_i;
 input [31:0] load_data_i;
 input [31:0] reset_adr_i;
 output [31:0] store_data_o;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire \u_decod.branch_imm_q_o[0] ;
 wire \u_decod.branch_imm_q_o[10] ;
 wire \u_decod.branch_imm_q_o[11] ;
 wire \u_decod.branch_imm_q_o[12] ;
 wire \u_decod.branch_imm_q_o[13] ;
 wire \u_decod.branch_imm_q_o[14] ;
 wire \u_decod.branch_imm_q_o[15] ;
 wire \u_decod.branch_imm_q_o[16] ;
 wire \u_decod.branch_imm_q_o[17] ;
 wire \u_decod.branch_imm_q_o[18] ;
 wire \u_decod.branch_imm_q_o[19] ;
 wire \u_decod.branch_imm_q_o[1] ;
 wire \u_decod.branch_imm_q_o[20] ;
 wire \u_decod.branch_imm_q_o[21] ;
 wire \u_decod.branch_imm_q_o[22] ;
 wire \u_decod.branch_imm_q_o[23] ;
 wire \u_decod.branch_imm_q_o[24] ;
 wire \u_decod.branch_imm_q_o[25] ;
 wire \u_decod.branch_imm_q_o[26] ;
 wire \u_decod.branch_imm_q_o[27] ;
 wire \u_decod.branch_imm_q_o[28] ;
 wire \u_decod.branch_imm_q_o[29] ;
 wire \u_decod.branch_imm_q_o[2] ;
 wire \u_decod.branch_imm_q_o[30] ;
 wire \u_decod.branch_imm_q_o[31] ;
 wire \u_decod.branch_imm_q_o[3] ;
 wire \u_decod.branch_imm_q_o[4] ;
 wire \u_decod.branch_imm_q_o[5] ;
 wire \u_decod.branch_imm_q_o[6] ;
 wire \u_decod.branch_imm_q_o[7] ;
 wire \u_decod.branch_imm_q_o[8] ;
 wire \u_decod.branch_imm_q_o[9] ;
 wire \u_decod.dec0.access_size_o[0] ;
 wire \u_decod.dec0.access_size_o[1] ;
 wire \u_decod.dec0.access_size_o[2] ;
 wire \u_decod.dec0.funct3[0] ;
 wire \u_decod.dec0.funct3[1] ;
 wire \u_decod.dec0.funct3[2] ;
 wire \u_decod.dec0.funct7[0] ;
 wire \u_decod.dec0.funct7[1] ;
 wire \u_decod.dec0.funct7[2] ;
 wire \u_decod.dec0.funct7[3] ;
 wire \u_decod.dec0.funct7[4] ;
 wire \u_decod.dec0.funct7[5] ;
 wire \u_decod.dec0.funct7[6] ;
 wire \u_decod.dec0.instr_i[0] ;
 wire \u_decod.dec0.instr_i[10] ;
 wire \u_decod.dec0.instr_i[11] ;
 wire \u_decod.dec0.instr_i[15] ;
 wire \u_decod.dec0.instr_i[16] ;
 wire \u_decod.dec0.instr_i[17] ;
 wire \u_decod.dec0.instr_i[18] ;
 wire \u_decod.dec0.instr_i[19] ;
 wire \u_decod.dec0.instr_i[1] ;
 wire \u_decod.dec0.instr_i[20] ;
 wire \u_decod.dec0.instr_i[21] ;
 wire \u_decod.dec0.instr_i[22] ;
 wire \u_decod.dec0.instr_i[23] ;
 wire \u_decod.dec0.instr_i[24] ;
 wire \u_decod.dec0.instr_i[2] ;
 wire \u_decod.dec0.instr_i[3] ;
 wire \u_decod.dec0.instr_i[4] ;
 wire \u_decod.dec0.instr_i[5] ;
 wire \u_decod.dec0.instr_i[6] ;
 wire \u_decod.dec0.instr_i[7] ;
 wire \u_decod.dec0.instr_i[8] ;
 wire \u_decod.dec0.instr_i[9] ;
 wire \u_decod.dec0.is_arithm ;
 wire \u_decod.dec0.is_branch ;
 wire \u_decod.dec0.is_shift ;
 wire \u_decod.dec0.jalr ;
 wire \u_decod.dec0.operation_o[0] ;
 wire \u_decod.dec0.operation_o[1] ;
 wire \u_decod.dec0.operation_o[2] ;
 wire \u_decod.dec0.operation_o[3] ;
 wire \u_decod.dec0.operation_o[4] ;
 wire \u_decod.dec0.rd_o[0] ;
 wire \u_decod.dec0.rd_o[1] ;
 wire \u_decod.dec0.rd_o[2] ;
 wire \u_decod.dec0.rd_o[3] ;
 wire \u_decod.dec0.rd_o[4] ;
 wire \u_decod.dec0.rd_v ;
 wire \u_decod.dec0.unit_o[3] ;
 wire \u_decod.dec0.unsign_extension ;
 wire \u_decod.exe_ff_rd_adr_q_i[0] ;
 wire \u_decod.exe_ff_rd_adr_q_i[1] ;
 wire \u_decod.exe_ff_rd_adr_q_i[2] ;
 wire \u_decod.exe_ff_rd_adr_q_i[3] ;
 wire \u_decod.exe_ff_rd_adr_q_i[4] ;
 wire \u_decod.exe_ff_res_data_i[0] ;
 wire \u_decod.exe_ff_res_data_i[10] ;
 wire \u_decod.exe_ff_res_data_i[11] ;
 wire \u_decod.exe_ff_res_data_i[12] ;
 wire \u_decod.exe_ff_res_data_i[13] ;
 wire \u_decod.exe_ff_res_data_i[14] ;
 wire \u_decod.exe_ff_res_data_i[15] ;
 wire \u_decod.exe_ff_res_data_i[16] ;
 wire \u_decod.exe_ff_res_data_i[17] ;
 wire \u_decod.exe_ff_res_data_i[18] ;
 wire \u_decod.exe_ff_res_data_i[19] ;
 wire \u_decod.exe_ff_res_data_i[1] ;
 wire \u_decod.exe_ff_res_data_i[20] ;
 wire \u_decod.exe_ff_res_data_i[21] ;
 wire \u_decod.exe_ff_res_data_i[22] ;
 wire \u_decod.exe_ff_res_data_i[23] ;
 wire \u_decod.exe_ff_res_data_i[24] ;
 wire \u_decod.exe_ff_res_data_i[25] ;
 wire \u_decod.exe_ff_res_data_i[26] ;
 wire \u_decod.exe_ff_res_data_i[27] ;
 wire \u_decod.exe_ff_res_data_i[28] ;
 wire \u_decod.exe_ff_res_data_i[29] ;
 wire \u_decod.exe_ff_res_data_i[2] ;
 wire \u_decod.exe_ff_res_data_i[30] ;
 wire \u_decod.exe_ff_res_data_i[31] ;
 wire \u_decod.exe_ff_res_data_i[3] ;
 wire \u_decod.exe_ff_res_data_i[4] ;
 wire \u_decod.exe_ff_res_data_i[5] ;
 wire \u_decod.exe_ff_res_data_i[6] ;
 wire \u_decod.exe_ff_res_data_i[7] ;
 wire \u_decod.exe_ff_res_data_i[8] ;
 wire \u_decod.exe_ff_res_data_i[9] ;
 wire \u_decod.exe_ff_write_v_q_i ;
 wire \u_decod.flush_v ;
 wire \u_decod.instr_operation_q[0] ;
 wire \u_decod.instr_operation_q[1] ;
 wire \u_decod.instr_operation_q[2] ;
 wire \u_decod.instr_operation_q[3] ;
 wire \u_decod.instr_operation_q[4] ;
 wire \u_decod.instr_operation_q[5] ;
 wire \u_decod.instr_unit_q[0] ;
 wire \u_decod.instr_unit_q[1] ;
 wire \u_decod.instr_unit_q[2] ;
 wire \u_decod.instr_unit_q[3] ;
 wire \u_decod.pc0_q_i[0] ;
 wire \u_decod.pc0_q_i[10] ;
 wire \u_decod.pc0_q_i[11] ;
 wire \u_decod.pc0_q_i[12] ;
 wire \u_decod.pc0_q_i[13] ;
 wire \u_decod.pc0_q_i[14] ;
 wire \u_decod.pc0_q_i[15] ;
 wire \u_decod.pc0_q_i[16] ;
 wire \u_decod.pc0_q_i[17] ;
 wire \u_decod.pc0_q_i[18] ;
 wire \u_decod.pc0_q_i[19] ;
 wire \u_decod.pc0_q_i[1] ;
 wire \u_decod.pc0_q_i[20] ;
 wire \u_decod.pc0_q_i[21] ;
 wire \u_decod.pc0_q_i[22] ;
 wire \u_decod.pc0_q_i[23] ;
 wire \u_decod.pc0_q_i[24] ;
 wire \u_decod.pc0_q_i[25] ;
 wire \u_decod.pc0_q_i[26] ;
 wire \u_decod.pc0_q_i[27] ;
 wire \u_decod.pc0_q_i[28] ;
 wire \u_decod.pc0_q_i[29] ;
 wire \u_decod.pc0_q_i[2] ;
 wire \u_decod.pc0_q_i[30] ;
 wire \u_decod.pc0_q_i[31] ;
 wire \u_decod.pc0_q_i[3] ;
 wire \u_decod.pc0_q_i[4] ;
 wire \u_decod.pc0_q_i[5] ;
 wire \u_decod.pc0_q_i[6] ;
 wire \u_decod.pc0_q_i[7] ;
 wire \u_decod.pc0_q_i[8] ;
 wire \u_decod.pc0_q_i[9] ;
 wire \u_decod.pc_q_o[0] ;
 wire \u_decod.pc_q_o[10] ;
 wire \u_decod.pc_q_o[11] ;
 wire \u_decod.pc_q_o[12] ;
 wire \u_decod.pc_q_o[13] ;
 wire \u_decod.pc_q_o[14] ;
 wire \u_decod.pc_q_o[15] ;
 wire \u_decod.pc_q_o[16] ;
 wire \u_decod.pc_q_o[17] ;
 wire \u_decod.pc_q_o[18] ;
 wire \u_decod.pc_q_o[19] ;
 wire \u_decod.pc_q_o[1] ;
 wire \u_decod.pc_q_o[20] ;
 wire \u_decod.pc_q_o[21] ;
 wire \u_decod.pc_q_o[22] ;
 wire \u_decod.pc_q_o[23] ;
 wire \u_decod.pc_q_o[24] ;
 wire \u_decod.pc_q_o[25] ;
 wire \u_decod.pc_q_o[26] ;
 wire \u_decod.pc_q_o[27] ;
 wire \u_decod.pc_q_o[28] ;
 wire \u_decod.pc_q_o[29] ;
 wire \u_decod.pc_q_o[2] ;
 wire \u_decod.pc_q_o[30] ;
 wire \u_decod.pc_q_o[31] ;
 wire \u_decod.pc_q_o[3] ;
 wire \u_decod.pc_q_o[4] ;
 wire \u_decod.pc_q_o[5] ;
 wire \u_decod.pc_q_o[6] ;
 wire \u_decod.pc_q_o[7] ;
 wire \u_decod.pc_q_o[8] ;
 wire \u_decod.pc_q_o[9] ;
 wire \u_decod.rd_v_q ;
 wire \u_decod.rf_ff_rd_adr_q_i[0] ;
 wire \u_decod.rf_ff_rd_adr_q_i[1] ;
 wire \u_decod.rf_ff_rd_adr_q_i[2] ;
 wire \u_decod.rf_ff_rd_adr_q_i[3] ;
 wire \u_decod.rf_ff_rd_adr_q_i[4] ;
 wire \u_decod.rf_ff_res_data_i[0] ;
 wire \u_decod.rf_ff_res_data_i[10] ;
 wire \u_decod.rf_ff_res_data_i[11] ;
 wire \u_decod.rf_ff_res_data_i[12] ;
 wire \u_decod.rf_ff_res_data_i[13] ;
 wire \u_decod.rf_ff_res_data_i[14] ;
 wire \u_decod.rf_ff_res_data_i[15] ;
 wire \u_decod.rf_ff_res_data_i[16] ;
 wire \u_decod.rf_ff_res_data_i[17] ;
 wire \u_decod.rf_ff_res_data_i[18] ;
 wire \u_decod.rf_ff_res_data_i[19] ;
 wire \u_decod.rf_ff_res_data_i[1] ;
 wire \u_decod.rf_ff_res_data_i[20] ;
 wire \u_decod.rf_ff_res_data_i[21] ;
 wire \u_decod.rf_ff_res_data_i[22] ;
 wire \u_decod.rf_ff_res_data_i[23] ;
 wire \u_decod.rf_ff_res_data_i[24] ;
 wire \u_decod.rf_ff_res_data_i[25] ;
 wire \u_decod.rf_ff_res_data_i[26] ;
 wire \u_decod.rf_ff_res_data_i[27] ;
 wire \u_decod.rf_ff_res_data_i[28] ;
 wire \u_decod.rf_ff_res_data_i[29] ;
 wire \u_decod.rf_ff_res_data_i[2] ;
 wire \u_decod.rf_ff_res_data_i[30] ;
 wire \u_decod.rf_ff_res_data_i[31] ;
 wire \u_decod.rf_ff_res_data_i[3] ;
 wire \u_decod.rf_ff_res_data_i[4] ;
 wire \u_decod.rf_ff_res_data_i[5] ;
 wire \u_decod.rf_ff_res_data_i[6] ;
 wire \u_decod.rf_ff_res_data_i[7] ;
 wire \u_decod.rf_ff_res_data_i[8] ;
 wire \u_decod.rf_ff_res_data_i[9] ;
 wire \u_decod.rf_write_v_q_i ;
 wire \u_decod.rs1_data[0] ;
 wire \u_decod.rs1_data[10] ;
 wire \u_decod.rs1_data[11] ;
 wire \u_decod.rs1_data[12] ;
 wire \u_decod.rs1_data[13] ;
 wire \u_decod.rs1_data[14] ;
 wire \u_decod.rs1_data[15] ;
 wire \u_decod.rs1_data[16] ;
 wire \u_decod.rs1_data[17] ;
 wire \u_decod.rs1_data[18] ;
 wire \u_decod.rs1_data[19] ;
 wire \u_decod.rs1_data[1] ;
 wire \u_decod.rs1_data[20] ;
 wire \u_decod.rs1_data[21] ;
 wire \u_decod.rs1_data[22] ;
 wire \u_decod.rs1_data[23] ;
 wire \u_decod.rs1_data[24] ;
 wire \u_decod.rs1_data[25] ;
 wire \u_decod.rs1_data[26] ;
 wire \u_decod.rs1_data[27] ;
 wire \u_decod.rs1_data[28] ;
 wire \u_decod.rs1_data[29] ;
 wire \u_decod.rs1_data[2] ;
 wire \u_decod.rs1_data[30] ;
 wire \u_decod.rs1_data[31] ;
 wire \u_decod.rs1_data[3] ;
 wire \u_decod.rs1_data[4] ;
 wire \u_decod.rs1_data[5] ;
 wire \u_decod.rs1_data[6] ;
 wire \u_decod.rs1_data[7] ;
 wire \u_decod.rs1_data[8] ;
 wire \u_decod.rs1_data[9] ;
 wire \u_decod.rs1_data_nxt[32] ;
 wire \u_decod.rs1_data_q[0] ;
 wire \u_decod.rs1_data_q[10] ;
 wire \u_decod.rs1_data_q[11] ;
 wire \u_decod.rs1_data_q[12] ;
 wire \u_decod.rs1_data_q[13] ;
 wire \u_decod.rs1_data_q[14] ;
 wire \u_decod.rs1_data_q[15] ;
 wire \u_decod.rs1_data_q[16] ;
 wire \u_decod.rs1_data_q[17] ;
 wire \u_decod.rs1_data_q[18] ;
 wire \u_decod.rs1_data_q[19] ;
 wire \u_decod.rs1_data_q[1] ;
 wire \u_decod.rs1_data_q[20] ;
 wire \u_decod.rs1_data_q[21] ;
 wire \u_decod.rs1_data_q[22] ;
 wire \u_decod.rs1_data_q[23] ;
 wire \u_decod.rs1_data_q[24] ;
 wire \u_decod.rs1_data_q[25] ;
 wire \u_decod.rs1_data_q[26] ;
 wire \u_decod.rs1_data_q[27] ;
 wire \u_decod.rs1_data_q[28] ;
 wire \u_decod.rs1_data_q[29] ;
 wire \u_decod.rs1_data_q[2] ;
 wire \u_decod.rs1_data_q[30] ;
 wire \u_decod.rs1_data_q[31] ;
 wire \u_decod.rs1_data_q[32] ;
 wire \u_decod.rs1_data_q[3] ;
 wire \u_decod.rs1_data_q[4] ;
 wire \u_decod.rs1_data_q[5] ;
 wire \u_decod.rs1_data_q[6] ;
 wire \u_decod.rs1_data_q[7] ;
 wire \u_decod.rs1_data_q[8] ;
 wire \u_decod.rs1_data_q[9] ;
 wire \u_decod.rs2_data_nxt[0] ;
 wire \u_decod.rs2_data_nxt[10] ;
 wire \u_decod.rs2_data_nxt[11] ;
 wire \u_decod.rs2_data_nxt[12] ;
 wire \u_decod.rs2_data_nxt[13] ;
 wire \u_decod.rs2_data_nxt[14] ;
 wire \u_decod.rs2_data_nxt[15] ;
 wire \u_decod.rs2_data_nxt[16] ;
 wire \u_decod.rs2_data_nxt[17] ;
 wire \u_decod.rs2_data_nxt[18] ;
 wire \u_decod.rs2_data_nxt[19] ;
 wire \u_decod.rs2_data_nxt[1] ;
 wire \u_decod.rs2_data_nxt[20] ;
 wire \u_decod.rs2_data_nxt[21] ;
 wire \u_decod.rs2_data_nxt[22] ;
 wire \u_decod.rs2_data_nxt[23] ;
 wire \u_decod.rs2_data_nxt[24] ;
 wire \u_decod.rs2_data_nxt[25] ;
 wire \u_decod.rs2_data_nxt[26] ;
 wire \u_decod.rs2_data_nxt[27] ;
 wire \u_decod.rs2_data_nxt[28] ;
 wire \u_decod.rs2_data_nxt[29] ;
 wire \u_decod.rs2_data_nxt[2] ;
 wire \u_decod.rs2_data_nxt[30] ;
 wire \u_decod.rs2_data_nxt[31] ;
 wire \u_decod.rs2_data_nxt[32] ;
 wire \u_decod.rs2_data_nxt[3] ;
 wire \u_decod.rs2_data_nxt[4] ;
 wire \u_decod.rs2_data_nxt[5] ;
 wire \u_decod.rs2_data_nxt[6] ;
 wire \u_decod.rs2_data_nxt[7] ;
 wire \u_decod.rs2_data_nxt[8] ;
 wire \u_decod.rs2_data_nxt[9] ;
 wire \u_decod.rs2_data_q[0] ;
 wire \u_decod.rs2_data_q[10] ;
 wire \u_decod.rs2_data_q[11] ;
 wire \u_decod.rs2_data_q[12] ;
 wire \u_decod.rs2_data_q[13] ;
 wire \u_decod.rs2_data_q[14] ;
 wire \u_decod.rs2_data_q[15] ;
 wire \u_decod.rs2_data_q[16] ;
 wire \u_decod.rs2_data_q[17] ;
 wire \u_decod.rs2_data_q[18] ;
 wire \u_decod.rs2_data_q[19] ;
 wire \u_decod.rs2_data_q[1] ;
 wire \u_decod.rs2_data_q[20] ;
 wire \u_decod.rs2_data_q[21] ;
 wire \u_decod.rs2_data_q[22] ;
 wire \u_decod.rs2_data_q[23] ;
 wire \u_decod.rs2_data_q[24] ;
 wire \u_decod.rs2_data_q[25] ;
 wire \u_decod.rs2_data_q[26] ;
 wire \u_decod.rs2_data_q[27] ;
 wire \u_decod.rs2_data_q[28] ;
 wire \u_decod.rs2_data_q[29] ;
 wire \u_decod.rs2_data_q[2] ;
 wire \u_decod.rs2_data_q[30] ;
 wire \u_decod.rs2_data_q[31] ;
 wire \u_decod.rs2_data_q[32] ;
 wire \u_decod.rs2_data_q[3] ;
 wire \u_decod.rs2_data_q[4] ;
 wire \u_decod.rs2_data_q[5] ;
 wire \u_decod.rs2_data_q[6] ;
 wire \u_decod.rs2_data_q[7] ;
 wire \u_decod.rs2_data_q[8] ;
 wire \u_decod.rs2_data_q[9] ;
 wire \u_decod.unsign_ext_q_o ;
 wire \u_exe.branch_v ;
 wire \u_exe.bu_pc_res[0] ;
 wire \u_exe.bu_pc_res[10] ;
 wire \u_exe.bu_pc_res[11] ;
 wire \u_exe.bu_pc_res[12] ;
 wire \u_exe.bu_pc_res[13] ;
 wire \u_exe.bu_pc_res[14] ;
 wire \u_exe.bu_pc_res[15] ;
 wire \u_exe.bu_pc_res[16] ;
 wire \u_exe.bu_pc_res[17] ;
 wire \u_exe.bu_pc_res[18] ;
 wire \u_exe.bu_pc_res[19] ;
 wire \u_exe.bu_pc_res[1] ;
 wire \u_exe.bu_pc_res[20] ;
 wire \u_exe.bu_pc_res[21] ;
 wire \u_exe.bu_pc_res[22] ;
 wire \u_exe.bu_pc_res[23] ;
 wire \u_exe.bu_pc_res[24] ;
 wire \u_exe.bu_pc_res[25] ;
 wire \u_exe.bu_pc_res[26] ;
 wire \u_exe.bu_pc_res[27] ;
 wire \u_exe.bu_pc_res[28] ;
 wire \u_exe.bu_pc_res[29] ;
 wire \u_exe.bu_pc_res[2] ;
 wire \u_exe.bu_pc_res[30] ;
 wire \u_exe.bu_pc_res[31] ;
 wire \u_exe.bu_pc_res[3] ;
 wire \u_exe.bu_pc_res[4] ;
 wire \u_exe.bu_pc_res[5] ;
 wire \u_exe.bu_pc_res[6] ;
 wire \u_exe.bu_pc_res[7] ;
 wire \u_exe.bu_pc_res[8] ;
 wire \u_exe.bu_pc_res[9] ;
 wire \u_exe.flush_v_dly1_q ;
 wire \u_exe.pc_data_q[0] ;
 wire \u_exe.pc_data_q[10] ;
 wire \u_exe.pc_data_q[11] ;
 wire \u_exe.pc_data_q[12] ;
 wire \u_exe.pc_data_q[13] ;
 wire \u_exe.pc_data_q[14] ;
 wire \u_exe.pc_data_q[15] ;
 wire \u_exe.pc_data_q[16] ;
 wire \u_exe.pc_data_q[17] ;
 wire \u_exe.pc_data_q[18] ;
 wire \u_exe.pc_data_q[19] ;
 wire \u_exe.pc_data_q[1] ;
 wire \u_exe.pc_data_q[20] ;
 wire \u_exe.pc_data_q[21] ;
 wire \u_exe.pc_data_q[22] ;
 wire \u_exe.pc_data_q[23] ;
 wire \u_exe.pc_data_q[24] ;
 wire \u_exe.pc_data_q[25] ;
 wire \u_exe.pc_data_q[26] ;
 wire \u_exe.pc_data_q[27] ;
 wire \u_exe.pc_data_q[28] ;
 wire \u_exe.pc_data_q[29] ;
 wire \u_exe.pc_data_q[2] ;
 wire \u_exe.pc_data_q[30] ;
 wire \u_exe.pc_data_q[31] ;
 wire \u_exe.pc_data_q[3] ;
 wire \u_exe.pc_data_q[4] ;
 wire \u_exe.pc_data_q[5] ;
 wire \u_exe.pc_data_q[6] ;
 wire \u_exe.pc_data_q[7] ;
 wire \u_exe.pc_data_q[8] ;
 wire \u_exe.pc_data_q[9] ;
 wire \u_ifetch.reset_n_q ;
 wire \u_rf.reg0_q[0] ;
 wire \u_rf.reg0_q[10] ;
 wire \u_rf.reg0_q[11] ;
 wire \u_rf.reg0_q[12] ;
 wire \u_rf.reg0_q[13] ;
 wire \u_rf.reg0_q[14] ;
 wire \u_rf.reg0_q[15] ;
 wire \u_rf.reg0_q[16] ;
 wire \u_rf.reg0_q[17] ;
 wire \u_rf.reg0_q[18] ;
 wire \u_rf.reg0_q[19] ;
 wire \u_rf.reg0_q[1] ;
 wire \u_rf.reg0_q[20] ;
 wire \u_rf.reg0_q[21] ;
 wire \u_rf.reg0_q[22] ;
 wire \u_rf.reg0_q[23] ;
 wire \u_rf.reg0_q[24] ;
 wire \u_rf.reg0_q[25] ;
 wire \u_rf.reg0_q[26] ;
 wire \u_rf.reg0_q[27] ;
 wire \u_rf.reg0_q[28] ;
 wire \u_rf.reg0_q[29] ;
 wire \u_rf.reg0_q[2] ;
 wire \u_rf.reg0_q[30] ;
 wire \u_rf.reg0_q[31] ;
 wire \u_rf.reg0_q[3] ;
 wire \u_rf.reg0_q[4] ;
 wire \u_rf.reg0_q[5] ;
 wire \u_rf.reg0_q[6] ;
 wire \u_rf.reg0_q[7] ;
 wire \u_rf.reg0_q[8] ;
 wire \u_rf.reg0_q[9] ;
 wire \u_rf.reg10_q[0] ;
 wire \u_rf.reg10_q[10] ;
 wire \u_rf.reg10_q[11] ;
 wire \u_rf.reg10_q[12] ;
 wire \u_rf.reg10_q[13] ;
 wire \u_rf.reg10_q[14] ;
 wire \u_rf.reg10_q[15] ;
 wire \u_rf.reg10_q[16] ;
 wire \u_rf.reg10_q[17] ;
 wire \u_rf.reg10_q[18] ;
 wire \u_rf.reg10_q[19] ;
 wire \u_rf.reg10_q[1] ;
 wire \u_rf.reg10_q[20] ;
 wire \u_rf.reg10_q[21] ;
 wire \u_rf.reg10_q[22] ;
 wire \u_rf.reg10_q[23] ;
 wire \u_rf.reg10_q[24] ;
 wire \u_rf.reg10_q[25] ;
 wire \u_rf.reg10_q[26] ;
 wire \u_rf.reg10_q[27] ;
 wire \u_rf.reg10_q[28] ;
 wire \u_rf.reg10_q[29] ;
 wire \u_rf.reg10_q[2] ;
 wire \u_rf.reg10_q[30] ;
 wire \u_rf.reg10_q[31] ;
 wire \u_rf.reg10_q[3] ;
 wire \u_rf.reg10_q[4] ;
 wire \u_rf.reg10_q[5] ;
 wire \u_rf.reg10_q[6] ;
 wire \u_rf.reg10_q[7] ;
 wire \u_rf.reg10_q[8] ;
 wire \u_rf.reg10_q[9] ;
 wire \u_rf.reg11_q[0] ;
 wire \u_rf.reg11_q[10] ;
 wire \u_rf.reg11_q[11] ;
 wire \u_rf.reg11_q[12] ;
 wire \u_rf.reg11_q[13] ;
 wire \u_rf.reg11_q[14] ;
 wire \u_rf.reg11_q[15] ;
 wire \u_rf.reg11_q[16] ;
 wire \u_rf.reg11_q[17] ;
 wire \u_rf.reg11_q[18] ;
 wire \u_rf.reg11_q[19] ;
 wire \u_rf.reg11_q[1] ;
 wire \u_rf.reg11_q[20] ;
 wire \u_rf.reg11_q[21] ;
 wire \u_rf.reg11_q[22] ;
 wire \u_rf.reg11_q[23] ;
 wire \u_rf.reg11_q[24] ;
 wire \u_rf.reg11_q[25] ;
 wire \u_rf.reg11_q[26] ;
 wire \u_rf.reg11_q[27] ;
 wire \u_rf.reg11_q[28] ;
 wire \u_rf.reg11_q[29] ;
 wire \u_rf.reg11_q[2] ;
 wire \u_rf.reg11_q[30] ;
 wire \u_rf.reg11_q[31] ;
 wire \u_rf.reg11_q[3] ;
 wire \u_rf.reg11_q[4] ;
 wire \u_rf.reg11_q[5] ;
 wire \u_rf.reg11_q[6] ;
 wire \u_rf.reg11_q[7] ;
 wire \u_rf.reg11_q[8] ;
 wire \u_rf.reg11_q[9] ;
 wire \u_rf.reg12_q[0] ;
 wire \u_rf.reg12_q[10] ;
 wire \u_rf.reg12_q[11] ;
 wire \u_rf.reg12_q[12] ;
 wire \u_rf.reg12_q[13] ;
 wire \u_rf.reg12_q[14] ;
 wire \u_rf.reg12_q[15] ;
 wire \u_rf.reg12_q[16] ;
 wire \u_rf.reg12_q[17] ;
 wire \u_rf.reg12_q[18] ;
 wire \u_rf.reg12_q[19] ;
 wire \u_rf.reg12_q[1] ;
 wire \u_rf.reg12_q[20] ;
 wire \u_rf.reg12_q[21] ;
 wire \u_rf.reg12_q[22] ;
 wire \u_rf.reg12_q[23] ;
 wire \u_rf.reg12_q[24] ;
 wire \u_rf.reg12_q[25] ;
 wire \u_rf.reg12_q[26] ;
 wire \u_rf.reg12_q[27] ;
 wire \u_rf.reg12_q[28] ;
 wire \u_rf.reg12_q[29] ;
 wire \u_rf.reg12_q[2] ;
 wire \u_rf.reg12_q[30] ;
 wire \u_rf.reg12_q[31] ;
 wire \u_rf.reg12_q[3] ;
 wire \u_rf.reg12_q[4] ;
 wire \u_rf.reg12_q[5] ;
 wire \u_rf.reg12_q[6] ;
 wire \u_rf.reg12_q[7] ;
 wire \u_rf.reg12_q[8] ;
 wire \u_rf.reg12_q[9] ;
 wire \u_rf.reg13_q[0] ;
 wire \u_rf.reg13_q[10] ;
 wire \u_rf.reg13_q[11] ;
 wire \u_rf.reg13_q[12] ;
 wire \u_rf.reg13_q[13] ;
 wire \u_rf.reg13_q[14] ;
 wire \u_rf.reg13_q[15] ;
 wire \u_rf.reg13_q[16] ;
 wire \u_rf.reg13_q[17] ;
 wire \u_rf.reg13_q[18] ;
 wire \u_rf.reg13_q[19] ;
 wire \u_rf.reg13_q[1] ;
 wire \u_rf.reg13_q[20] ;
 wire \u_rf.reg13_q[21] ;
 wire \u_rf.reg13_q[22] ;
 wire \u_rf.reg13_q[23] ;
 wire \u_rf.reg13_q[24] ;
 wire \u_rf.reg13_q[25] ;
 wire \u_rf.reg13_q[26] ;
 wire \u_rf.reg13_q[27] ;
 wire \u_rf.reg13_q[28] ;
 wire \u_rf.reg13_q[29] ;
 wire \u_rf.reg13_q[2] ;
 wire \u_rf.reg13_q[30] ;
 wire \u_rf.reg13_q[31] ;
 wire \u_rf.reg13_q[3] ;
 wire \u_rf.reg13_q[4] ;
 wire \u_rf.reg13_q[5] ;
 wire \u_rf.reg13_q[6] ;
 wire \u_rf.reg13_q[7] ;
 wire \u_rf.reg13_q[8] ;
 wire \u_rf.reg13_q[9] ;
 wire \u_rf.reg14_q[0] ;
 wire \u_rf.reg14_q[10] ;
 wire \u_rf.reg14_q[11] ;
 wire \u_rf.reg14_q[12] ;
 wire \u_rf.reg14_q[13] ;
 wire \u_rf.reg14_q[14] ;
 wire \u_rf.reg14_q[15] ;
 wire \u_rf.reg14_q[16] ;
 wire \u_rf.reg14_q[17] ;
 wire \u_rf.reg14_q[18] ;
 wire \u_rf.reg14_q[19] ;
 wire \u_rf.reg14_q[1] ;
 wire \u_rf.reg14_q[20] ;
 wire \u_rf.reg14_q[21] ;
 wire \u_rf.reg14_q[22] ;
 wire \u_rf.reg14_q[23] ;
 wire \u_rf.reg14_q[24] ;
 wire \u_rf.reg14_q[25] ;
 wire \u_rf.reg14_q[26] ;
 wire \u_rf.reg14_q[27] ;
 wire \u_rf.reg14_q[28] ;
 wire \u_rf.reg14_q[29] ;
 wire \u_rf.reg14_q[2] ;
 wire \u_rf.reg14_q[30] ;
 wire \u_rf.reg14_q[31] ;
 wire \u_rf.reg14_q[3] ;
 wire \u_rf.reg14_q[4] ;
 wire \u_rf.reg14_q[5] ;
 wire \u_rf.reg14_q[6] ;
 wire \u_rf.reg14_q[7] ;
 wire \u_rf.reg14_q[8] ;
 wire \u_rf.reg14_q[9] ;
 wire \u_rf.reg15_q[0] ;
 wire \u_rf.reg15_q[10] ;
 wire \u_rf.reg15_q[11] ;
 wire \u_rf.reg15_q[12] ;
 wire \u_rf.reg15_q[13] ;
 wire \u_rf.reg15_q[14] ;
 wire \u_rf.reg15_q[15] ;
 wire \u_rf.reg15_q[16] ;
 wire \u_rf.reg15_q[17] ;
 wire \u_rf.reg15_q[18] ;
 wire \u_rf.reg15_q[19] ;
 wire \u_rf.reg15_q[1] ;
 wire \u_rf.reg15_q[20] ;
 wire \u_rf.reg15_q[21] ;
 wire \u_rf.reg15_q[22] ;
 wire \u_rf.reg15_q[23] ;
 wire \u_rf.reg15_q[24] ;
 wire \u_rf.reg15_q[25] ;
 wire \u_rf.reg15_q[26] ;
 wire \u_rf.reg15_q[27] ;
 wire \u_rf.reg15_q[28] ;
 wire \u_rf.reg15_q[29] ;
 wire \u_rf.reg15_q[2] ;
 wire \u_rf.reg15_q[30] ;
 wire \u_rf.reg15_q[31] ;
 wire \u_rf.reg15_q[3] ;
 wire \u_rf.reg15_q[4] ;
 wire \u_rf.reg15_q[5] ;
 wire \u_rf.reg15_q[6] ;
 wire \u_rf.reg15_q[7] ;
 wire \u_rf.reg15_q[8] ;
 wire \u_rf.reg15_q[9] ;
 wire \u_rf.reg16_q[0] ;
 wire \u_rf.reg16_q[10] ;
 wire \u_rf.reg16_q[11] ;
 wire \u_rf.reg16_q[12] ;
 wire \u_rf.reg16_q[13] ;
 wire \u_rf.reg16_q[14] ;
 wire \u_rf.reg16_q[15] ;
 wire \u_rf.reg16_q[16] ;
 wire \u_rf.reg16_q[17] ;
 wire \u_rf.reg16_q[18] ;
 wire \u_rf.reg16_q[19] ;
 wire \u_rf.reg16_q[1] ;
 wire \u_rf.reg16_q[20] ;
 wire \u_rf.reg16_q[21] ;
 wire \u_rf.reg16_q[22] ;
 wire \u_rf.reg16_q[23] ;
 wire \u_rf.reg16_q[24] ;
 wire \u_rf.reg16_q[25] ;
 wire \u_rf.reg16_q[26] ;
 wire \u_rf.reg16_q[27] ;
 wire \u_rf.reg16_q[28] ;
 wire \u_rf.reg16_q[29] ;
 wire \u_rf.reg16_q[2] ;
 wire \u_rf.reg16_q[30] ;
 wire \u_rf.reg16_q[31] ;
 wire \u_rf.reg16_q[3] ;
 wire \u_rf.reg16_q[4] ;
 wire \u_rf.reg16_q[5] ;
 wire \u_rf.reg16_q[6] ;
 wire \u_rf.reg16_q[7] ;
 wire \u_rf.reg16_q[8] ;
 wire \u_rf.reg16_q[9] ;
 wire \u_rf.reg17_q[0] ;
 wire \u_rf.reg17_q[10] ;
 wire \u_rf.reg17_q[11] ;
 wire \u_rf.reg17_q[12] ;
 wire \u_rf.reg17_q[13] ;
 wire \u_rf.reg17_q[14] ;
 wire \u_rf.reg17_q[15] ;
 wire \u_rf.reg17_q[16] ;
 wire \u_rf.reg17_q[17] ;
 wire \u_rf.reg17_q[18] ;
 wire \u_rf.reg17_q[19] ;
 wire \u_rf.reg17_q[1] ;
 wire \u_rf.reg17_q[20] ;
 wire \u_rf.reg17_q[21] ;
 wire \u_rf.reg17_q[22] ;
 wire \u_rf.reg17_q[23] ;
 wire \u_rf.reg17_q[24] ;
 wire \u_rf.reg17_q[25] ;
 wire \u_rf.reg17_q[26] ;
 wire \u_rf.reg17_q[27] ;
 wire \u_rf.reg17_q[28] ;
 wire \u_rf.reg17_q[29] ;
 wire \u_rf.reg17_q[2] ;
 wire \u_rf.reg17_q[30] ;
 wire \u_rf.reg17_q[31] ;
 wire \u_rf.reg17_q[3] ;
 wire \u_rf.reg17_q[4] ;
 wire \u_rf.reg17_q[5] ;
 wire \u_rf.reg17_q[6] ;
 wire \u_rf.reg17_q[7] ;
 wire \u_rf.reg17_q[8] ;
 wire \u_rf.reg17_q[9] ;
 wire \u_rf.reg18_q[0] ;
 wire \u_rf.reg18_q[10] ;
 wire \u_rf.reg18_q[11] ;
 wire \u_rf.reg18_q[12] ;
 wire \u_rf.reg18_q[13] ;
 wire \u_rf.reg18_q[14] ;
 wire \u_rf.reg18_q[15] ;
 wire \u_rf.reg18_q[16] ;
 wire \u_rf.reg18_q[17] ;
 wire \u_rf.reg18_q[18] ;
 wire \u_rf.reg18_q[19] ;
 wire \u_rf.reg18_q[1] ;
 wire \u_rf.reg18_q[20] ;
 wire \u_rf.reg18_q[21] ;
 wire \u_rf.reg18_q[22] ;
 wire \u_rf.reg18_q[23] ;
 wire \u_rf.reg18_q[24] ;
 wire \u_rf.reg18_q[25] ;
 wire \u_rf.reg18_q[26] ;
 wire \u_rf.reg18_q[27] ;
 wire \u_rf.reg18_q[28] ;
 wire \u_rf.reg18_q[29] ;
 wire \u_rf.reg18_q[2] ;
 wire \u_rf.reg18_q[30] ;
 wire \u_rf.reg18_q[31] ;
 wire \u_rf.reg18_q[3] ;
 wire \u_rf.reg18_q[4] ;
 wire \u_rf.reg18_q[5] ;
 wire \u_rf.reg18_q[6] ;
 wire \u_rf.reg18_q[7] ;
 wire \u_rf.reg18_q[8] ;
 wire \u_rf.reg18_q[9] ;
 wire \u_rf.reg19_q[0] ;
 wire \u_rf.reg19_q[10] ;
 wire \u_rf.reg19_q[11] ;
 wire \u_rf.reg19_q[12] ;
 wire \u_rf.reg19_q[13] ;
 wire \u_rf.reg19_q[14] ;
 wire \u_rf.reg19_q[15] ;
 wire \u_rf.reg19_q[16] ;
 wire \u_rf.reg19_q[17] ;
 wire \u_rf.reg19_q[18] ;
 wire \u_rf.reg19_q[19] ;
 wire \u_rf.reg19_q[1] ;
 wire \u_rf.reg19_q[20] ;
 wire \u_rf.reg19_q[21] ;
 wire \u_rf.reg19_q[22] ;
 wire \u_rf.reg19_q[23] ;
 wire \u_rf.reg19_q[24] ;
 wire \u_rf.reg19_q[25] ;
 wire \u_rf.reg19_q[26] ;
 wire \u_rf.reg19_q[27] ;
 wire \u_rf.reg19_q[28] ;
 wire \u_rf.reg19_q[29] ;
 wire \u_rf.reg19_q[2] ;
 wire \u_rf.reg19_q[30] ;
 wire \u_rf.reg19_q[31] ;
 wire \u_rf.reg19_q[3] ;
 wire \u_rf.reg19_q[4] ;
 wire \u_rf.reg19_q[5] ;
 wire \u_rf.reg19_q[6] ;
 wire \u_rf.reg19_q[7] ;
 wire \u_rf.reg19_q[8] ;
 wire \u_rf.reg19_q[9] ;
 wire \u_rf.reg1_q[0] ;
 wire \u_rf.reg1_q[10] ;
 wire \u_rf.reg1_q[11] ;
 wire \u_rf.reg1_q[12] ;
 wire \u_rf.reg1_q[13] ;
 wire \u_rf.reg1_q[14] ;
 wire \u_rf.reg1_q[15] ;
 wire \u_rf.reg1_q[16] ;
 wire \u_rf.reg1_q[17] ;
 wire \u_rf.reg1_q[18] ;
 wire \u_rf.reg1_q[19] ;
 wire \u_rf.reg1_q[1] ;
 wire \u_rf.reg1_q[20] ;
 wire \u_rf.reg1_q[21] ;
 wire \u_rf.reg1_q[22] ;
 wire \u_rf.reg1_q[23] ;
 wire \u_rf.reg1_q[24] ;
 wire \u_rf.reg1_q[25] ;
 wire \u_rf.reg1_q[26] ;
 wire \u_rf.reg1_q[27] ;
 wire \u_rf.reg1_q[28] ;
 wire \u_rf.reg1_q[29] ;
 wire \u_rf.reg1_q[2] ;
 wire \u_rf.reg1_q[30] ;
 wire \u_rf.reg1_q[31] ;
 wire \u_rf.reg1_q[3] ;
 wire \u_rf.reg1_q[4] ;
 wire \u_rf.reg1_q[5] ;
 wire \u_rf.reg1_q[6] ;
 wire \u_rf.reg1_q[7] ;
 wire \u_rf.reg1_q[8] ;
 wire \u_rf.reg1_q[9] ;
 wire \u_rf.reg20_q[0] ;
 wire \u_rf.reg20_q[10] ;
 wire \u_rf.reg20_q[11] ;
 wire \u_rf.reg20_q[12] ;
 wire \u_rf.reg20_q[13] ;
 wire \u_rf.reg20_q[14] ;
 wire \u_rf.reg20_q[15] ;
 wire \u_rf.reg20_q[16] ;
 wire \u_rf.reg20_q[17] ;
 wire \u_rf.reg20_q[18] ;
 wire \u_rf.reg20_q[19] ;
 wire \u_rf.reg20_q[1] ;
 wire \u_rf.reg20_q[20] ;
 wire \u_rf.reg20_q[21] ;
 wire \u_rf.reg20_q[22] ;
 wire \u_rf.reg20_q[23] ;
 wire \u_rf.reg20_q[24] ;
 wire \u_rf.reg20_q[25] ;
 wire \u_rf.reg20_q[26] ;
 wire \u_rf.reg20_q[27] ;
 wire \u_rf.reg20_q[28] ;
 wire \u_rf.reg20_q[29] ;
 wire \u_rf.reg20_q[2] ;
 wire \u_rf.reg20_q[30] ;
 wire \u_rf.reg20_q[31] ;
 wire \u_rf.reg20_q[3] ;
 wire \u_rf.reg20_q[4] ;
 wire \u_rf.reg20_q[5] ;
 wire \u_rf.reg20_q[6] ;
 wire \u_rf.reg20_q[7] ;
 wire \u_rf.reg20_q[8] ;
 wire \u_rf.reg20_q[9] ;
 wire \u_rf.reg21_q[0] ;
 wire \u_rf.reg21_q[10] ;
 wire \u_rf.reg21_q[11] ;
 wire \u_rf.reg21_q[12] ;
 wire \u_rf.reg21_q[13] ;
 wire \u_rf.reg21_q[14] ;
 wire \u_rf.reg21_q[15] ;
 wire \u_rf.reg21_q[16] ;
 wire \u_rf.reg21_q[17] ;
 wire \u_rf.reg21_q[18] ;
 wire \u_rf.reg21_q[19] ;
 wire \u_rf.reg21_q[1] ;
 wire \u_rf.reg21_q[20] ;
 wire \u_rf.reg21_q[21] ;
 wire \u_rf.reg21_q[22] ;
 wire \u_rf.reg21_q[23] ;
 wire \u_rf.reg21_q[24] ;
 wire \u_rf.reg21_q[25] ;
 wire \u_rf.reg21_q[26] ;
 wire \u_rf.reg21_q[27] ;
 wire \u_rf.reg21_q[28] ;
 wire \u_rf.reg21_q[29] ;
 wire \u_rf.reg21_q[2] ;
 wire \u_rf.reg21_q[30] ;
 wire \u_rf.reg21_q[31] ;
 wire \u_rf.reg21_q[3] ;
 wire \u_rf.reg21_q[4] ;
 wire \u_rf.reg21_q[5] ;
 wire \u_rf.reg21_q[6] ;
 wire \u_rf.reg21_q[7] ;
 wire \u_rf.reg21_q[8] ;
 wire \u_rf.reg21_q[9] ;
 wire \u_rf.reg22_q[0] ;
 wire \u_rf.reg22_q[10] ;
 wire \u_rf.reg22_q[11] ;
 wire \u_rf.reg22_q[12] ;
 wire \u_rf.reg22_q[13] ;
 wire \u_rf.reg22_q[14] ;
 wire \u_rf.reg22_q[15] ;
 wire \u_rf.reg22_q[16] ;
 wire \u_rf.reg22_q[17] ;
 wire \u_rf.reg22_q[18] ;
 wire \u_rf.reg22_q[19] ;
 wire \u_rf.reg22_q[1] ;
 wire \u_rf.reg22_q[20] ;
 wire \u_rf.reg22_q[21] ;
 wire \u_rf.reg22_q[22] ;
 wire \u_rf.reg22_q[23] ;
 wire \u_rf.reg22_q[24] ;
 wire \u_rf.reg22_q[25] ;
 wire \u_rf.reg22_q[26] ;
 wire \u_rf.reg22_q[27] ;
 wire \u_rf.reg22_q[28] ;
 wire \u_rf.reg22_q[29] ;
 wire \u_rf.reg22_q[2] ;
 wire \u_rf.reg22_q[30] ;
 wire \u_rf.reg22_q[31] ;
 wire \u_rf.reg22_q[3] ;
 wire \u_rf.reg22_q[4] ;
 wire \u_rf.reg22_q[5] ;
 wire \u_rf.reg22_q[6] ;
 wire \u_rf.reg22_q[7] ;
 wire \u_rf.reg22_q[8] ;
 wire \u_rf.reg22_q[9] ;
 wire \u_rf.reg23_q[0] ;
 wire \u_rf.reg23_q[10] ;
 wire \u_rf.reg23_q[11] ;
 wire \u_rf.reg23_q[12] ;
 wire \u_rf.reg23_q[13] ;
 wire \u_rf.reg23_q[14] ;
 wire \u_rf.reg23_q[15] ;
 wire \u_rf.reg23_q[16] ;
 wire \u_rf.reg23_q[17] ;
 wire \u_rf.reg23_q[18] ;
 wire \u_rf.reg23_q[19] ;
 wire \u_rf.reg23_q[1] ;
 wire \u_rf.reg23_q[20] ;
 wire \u_rf.reg23_q[21] ;
 wire \u_rf.reg23_q[22] ;
 wire \u_rf.reg23_q[23] ;
 wire \u_rf.reg23_q[24] ;
 wire \u_rf.reg23_q[25] ;
 wire \u_rf.reg23_q[26] ;
 wire \u_rf.reg23_q[27] ;
 wire \u_rf.reg23_q[28] ;
 wire \u_rf.reg23_q[29] ;
 wire \u_rf.reg23_q[2] ;
 wire \u_rf.reg23_q[30] ;
 wire \u_rf.reg23_q[31] ;
 wire \u_rf.reg23_q[3] ;
 wire \u_rf.reg23_q[4] ;
 wire \u_rf.reg23_q[5] ;
 wire \u_rf.reg23_q[6] ;
 wire \u_rf.reg23_q[7] ;
 wire \u_rf.reg23_q[8] ;
 wire \u_rf.reg23_q[9] ;
 wire \u_rf.reg24_q[0] ;
 wire \u_rf.reg24_q[10] ;
 wire \u_rf.reg24_q[11] ;
 wire \u_rf.reg24_q[12] ;
 wire \u_rf.reg24_q[13] ;
 wire \u_rf.reg24_q[14] ;
 wire \u_rf.reg24_q[15] ;
 wire \u_rf.reg24_q[16] ;
 wire \u_rf.reg24_q[17] ;
 wire \u_rf.reg24_q[18] ;
 wire \u_rf.reg24_q[19] ;
 wire \u_rf.reg24_q[1] ;
 wire \u_rf.reg24_q[20] ;
 wire \u_rf.reg24_q[21] ;
 wire \u_rf.reg24_q[22] ;
 wire \u_rf.reg24_q[23] ;
 wire \u_rf.reg24_q[24] ;
 wire \u_rf.reg24_q[25] ;
 wire \u_rf.reg24_q[26] ;
 wire \u_rf.reg24_q[27] ;
 wire \u_rf.reg24_q[28] ;
 wire \u_rf.reg24_q[29] ;
 wire \u_rf.reg24_q[2] ;
 wire \u_rf.reg24_q[30] ;
 wire \u_rf.reg24_q[31] ;
 wire \u_rf.reg24_q[3] ;
 wire \u_rf.reg24_q[4] ;
 wire \u_rf.reg24_q[5] ;
 wire \u_rf.reg24_q[6] ;
 wire \u_rf.reg24_q[7] ;
 wire \u_rf.reg24_q[8] ;
 wire \u_rf.reg24_q[9] ;
 wire \u_rf.reg25_q[0] ;
 wire \u_rf.reg25_q[10] ;
 wire \u_rf.reg25_q[11] ;
 wire \u_rf.reg25_q[12] ;
 wire \u_rf.reg25_q[13] ;
 wire \u_rf.reg25_q[14] ;
 wire \u_rf.reg25_q[15] ;
 wire \u_rf.reg25_q[16] ;
 wire \u_rf.reg25_q[17] ;
 wire \u_rf.reg25_q[18] ;
 wire \u_rf.reg25_q[19] ;
 wire \u_rf.reg25_q[1] ;
 wire \u_rf.reg25_q[20] ;
 wire \u_rf.reg25_q[21] ;
 wire \u_rf.reg25_q[22] ;
 wire \u_rf.reg25_q[23] ;
 wire \u_rf.reg25_q[24] ;
 wire \u_rf.reg25_q[25] ;
 wire \u_rf.reg25_q[26] ;
 wire \u_rf.reg25_q[27] ;
 wire \u_rf.reg25_q[28] ;
 wire \u_rf.reg25_q[29] ;
 wire \u_rf.reg25_q[2] ;
 wire \u_rf.reg25_q[30] ;
 wire \u_rf.reg25_q[31] ;
 wire \u_rf.reg25_q[3] ;
 wire \u_rf.reg25_q[4] ;
 wire \u_rf.reg25_q[5] ;
 wire \u_rf.reg25_q[6] ;
 wire \u_rf.reg25_q[7] ;
 wire \u_rf.reg25_q[8] ;
 wire \u_rf.reg25_q[9] ;
 wire \u_rf.reg26_q[0] ;
 wire \u_rf.reg26_q[10] ;
 wire \u_rf.reg26_q[11] ;
 wire \u_rf.reg26_q[12] ;
 wire \u_rf.reg26_q[13] ;
 wire \u_rf.reg26_q[14] ;
 wire \u_rf.reg26_q[15] ;
 wire \u_rf.reg26_q[16] ;
 wire \u_rf.reg26_q[17] ;
 wire \u_rf.reg26_q[18] ;
 wire \u_rf.reg26_q[19] ;
 wire \u_rf.reg26_q[1] ;
 wire \u_rf.reg26_q[20] ;
 wire \u_rf.reg26_q[21] ;
 wire \u_rf.reg26_q[22] ;
 wire \u_rf.reg26_q[23] ;
 wire \u_rf.reg26_q[24] ;
 wire \u_rf.reg26_q[25] ;
 wire \u_rf.reg26_q[26] ;
 wire \u_rf.reg26_q[27] ;
 wire \u_rf.reg26_q[28] ;
 wire \u_rf.reg26_q[29] ;
 wire \u_rf.reg26_q[2] ;
 wire \u_rf.reg26_q[30] ;
 wire \u_rf.reg26_q[31] ;
 wire \u_rf.reg26_q[3] ;
 wire \u_rf.reg26_q[4] ;
 wire \u_rf.reg26_q[5] ;
 wire \u_rf.reg26_q[6] ;
 wire \u_rf.reg26_q[7] ;
 wire \u_rf.reg26_q[8] ;
 wire \u_rf.reg26_q[9] ;
 wire \u_rf.reg27_q[0] ;
 wire \u_rf.reg27_q[10] ;
 wire \u_rf.reg27_q[11] ;
 wire \u_rf.reg27_q[12] ;
 wire \u_rf.reg27_q[13] ;
 wire \u_rf.reg27_q[14] ;
 wire \u_rf.reg27_q[15] ;
 wire \u_rf.reg27_q[16] ;
 wire \u_rf.reg27_q[17] ;
 wire \u_rf.reg27_q[18] ;
 wire \u_rf.reg27_q[19] ;
 wire \u_rf.reg27_q[1] ;
 wire \u_rf.reg27_q[20] ;
 wire \u_rf.reg27_q[21] ;
 wire \u_rf.reg27_q[22] ;
 wire \u_rf.reg27_q[23] ;
 wire \u_rf.reg27_q[24] ;
 wire \u_rf.reg27_q[25] ;
 wire \u_rf.reg27_q[26] ;
 wire \u_rf.reg27_q[27] ;
 wire \u_rf.reg27_q[28] ;
 wire \u_rf.reg27_q[29] ;
 wire \u_rf.reg27_q[2] ;
 wire \u_rf.reg27_q[30] ;
 wire \u_rf.reg27_q[31] ;
 wire \u_rf.reg27_q[3] ;
 wire \u_rf.reg27_q[4] ;
 wire \u_rf.reg27_q[5] ;
 wire \u_rf.reg27_q[6] ;
 wire \u_rf.reg27_q[7] ;
 wire \u_rf.reg27_q[8] ;
 wire \u_rf.reg27_q[9] ;
 wire \u_rf.reg28_q[0] ;
 wire \u_rf.reg28_q[10] ;
 wire \u_rf.reg28_q[11] ;
 wire \u_rf.reg28_q[12] ;
 wire \u_rf.reg28_q[13] ;
 wire \u_rf.reg28_q[14] ;
 wire \u_rf.reg28_q[15] ;
 wire \u_rf.reg28_q[16] ;
 wire \u_rf.reg28_q[17] ;
 wire \u_rf.reg28_q[18] ;
 wire \u_rf.reg28_q[19] ;
 wire \u_rf.reg28_q[1] ;
 wire \u_rf.reg28_q[20] ;
 wire \u_rf.reg28_q[21] ;
 wire \u_rf.reg28_q[22] ;
 wire \u_rf.reg28_q[23] ;
 wire \u_rf.reg28_q[24] ;
 wire \u_rf.reg28_q[25] ;
 wire \u_rf.reg28_q[26] ;
 wire \u_rf.reg28_q[27] ;
 wire \u_rf.reg28_q[28] ;
 wire \u_rf.reg28_q[29] ;
 wire \u_rf.reg28_q[2] ;
 wire \u_rf.reg28_q[30] ;
 wire \u_rf.reg28_q[31] ;
 wire \u_rf.reg28_q[3] ;
 wire \u_rf.reg28_q[4] ;
 wire \u_rf.reg28_q[5] ;
 wire \u_rf.reg28_q[6] ;
 wire \u_rf.reg28_q[7] ;
 wire \u_rf.reg28_q[8] ;
 wire \u_rf.reg28_q[9] ;
 wire \u_rf.reg29_q[0] ;
 wire \u_rf.reg29_q[10] ;
 wire \u_rf.reg29_q[11] ;
 wire \u_rf.reg29_q[12] ;
 wire \u_rf.reg29_q[13] ;
 wire \u_rf.reg29_q[14] ;
 wire \u_rf.reg29_q[15] ;
 wire \u_rf.reg29_q[16] ;
 wire \u_rf.reg29_q[17] ;
 wire \u_rf.reg29_q[18] ;
 wire \u_rf.reg29_q[19] ;
 wire \u_rf.reg29_q[1] ;
 wire \u_rf.reg29_q[20] ;
 wire \u_rf.reg29_q[21] ;
 wire \u_rf.reg29_q[22] ;
 wire \u_rf.reg29_q[23] ;
 wire \u_rf.reg29_q[24] ;
 wire \u_rf.reg29_q[25] ;
 wire \u_rf.reg29_q[26] ;
 wire \u_rf.reg29_q[27] ;
 wire \u_rf.reg29_q[28] ;
 wire \u_rf.reg29_q[29] ;
 wire \u_rf.reg29_q[2] ;
 wire \u_rf.reg29_q[30] ;
 wire \u_rf.reg29_q[31] ;
 wire \u_rf.reg29_q[3] ;
 wire \u_rf.reg29_q[4] ;
 wire \u_rf.reg29_q[5] ;
 wire \u_rf.reg29_q[6] ;
 wire \u_rf.reg29_q[7] ;
 wire \u_rf.reg29_q[8] ;
 wire \u_rf.reg29_q[9] ;
 wire \u_rf.reg2_q[0] ;
 wire \u_rf.reg2_q[10] ;
 wire \u_rf.reg2_q[11] ;
 wire \u_rf.reg2_q[12] ;
 wire \u_rf.reg2_q[13] ;
 wire \u_rf.reg2_q[14] ;
 wire \u_rf.reg2_q[15] ;
 wire \u_rf.reg2_q[16] ;
 wire \u_rf.reg2_q[17] ;
 wire \u_rf.reg2_q[18] ;
 wire \u_rf.reg2_q[19] ;
 wire \u_rf.reg2_q[1] ;
 wire \u_rf.reg2_q[20] ;
 wire \u_rf.reg2_q[21] ;
 wire \u_rf.reg2_q[22] ;
 wire \u_rf.reg2_q[23] ;
 wire \u_rf.reg2_q[24] ;
 wire \u_rf.reg2_q[25] ;
 wire \u_rf.reg2_q[26] ;
 wire \u_rf.reg2_q[27] ;
 wire \u_rf.reg2_q[28] ;
 wire \u_rf.reg2_q[29] ;
 wire \u_rf.reg2_q[2] ;
 wire \u_rf.reg2_q[30] ;
 wire \u_rf.reg2_q[31] ;
 wire \u_rf.reg2_q[3] ;
 wire \u_rf.reg2_q[4] ;
 wire \u_rf.reg2_q[5] ;
 wire \u_rf.reg2_q[6] ;
 wire \u_rf.reg2_q[7] ;
 wire \u_rf.reg2_q[8] ;
 wire \u_rf.reg2_q[9] ;
 wire \u_rf.reg30_q[0] ;
 wire \u_rf.reg30_q[10] ;
 wire \u_rf.reg30_q[11] ;
 wire \u_rf.reg30_q[12] ;
 wire \u_rf.reg30_q[13] ;
 wire \u_rf.reg30_q[14] ;
 wire \u_rf.reg30_q[15] ;
 wire \u_rf.reg30_q[16] ;
 wire \u_rf.reg30_q[17] ;
 wire \u_rf.reg30_q[18] ;
 wire \u_rf.reg30_q[19] ;
 wire \u_rf.reg30_q[1] ;
 wire \u_rf.reg30_q[20] ;
 wire \u_rf.reg30_q[21] ;
 wire \u_rf.reg30_q[22] ;
 wire \u_rf.reg30_q[23] ;
 wire \u_rf.reg30_q[24] ;
 wire \u_rf.reg30_q[25] ;
 wire \u_rf.reg30_q[26] ;
 wire \u_rf.reg30_q[27] ;
 wire \u_rf.reg30_q[28] ;
 wire \u_rf.reg30_q[29] ;
 wire \u_rf.reg30_q[2] ;
 wire \u_rf.reg30_q[30] ;
 wire \u_rf.reg30_q[31] ;
 wire \u_rf.reg30_q[3] ;
 wire \u_rf.reg30_q[4] ;
 wire \u_rf.reg30_q[5] ;
 wire \u_rf.reg30_q[6] ;
 wire \u_rf.reg30_q[7] ;
 wire \u_rf.reg30_q[8] ;
 wire \u_rf.reg30_q[9] ;
 wire \u_rf.reg31_q[0] ;
 wire \u_rf.reg31_q[10] ;
 wire \u_rf.reg31_q[11] ;
 wire \u_rf.reg31_q[12] ;
 wire \u_rf.reg31_q[13] ;
 wire \u_rf.reg31_q[14] ;
 wire \u_rf.reg31_q[15] ;
 wire \u_rf.reg31_q[16] ;
 wire \u_rf.reg31_q[17] ;
 wire \u_rf.reg31_q[18] ;
 wire \u_rf.reg31_q[19] ;
 wire \u_rf.reg31_q[1] ;
 wire \u_rf.reg31_q[20] ;
 wire \u_rf.reg31_q[21] ;
 wire \u_rf.reg31_q[22] ;
 wire \u_rf.reg31_q[23] ;
 wire \u_rf.reg31_q[24] ;
 wire \u_rf.reg31_q[25] ;
 wire \u_rf.reg31_q[26] ;
 wire \u_rf.reg31_q[27] ;
 wire \u_rf.reg31_q[28] ;
 wire \u_rf.reg31_q[29] ;
 wire \u_rf.reg31_q[2] ;
 wire \u_rf.reg31_q[30] ;
 wire \u_rf.reg31_q[31] ;
 wire \u_rf.reg31_q[3] ;
 wire \u_rf.reg31_q[4] ;
 wire \u_rf.reg31_q[5] ;
 wire \u_rf.reg31_q[6] ;
 wire \u_rf.reg31_q[7] ;
 wire \u_rf.reg31_q[8] ;
 wire \u_rf.reg31_q[9] ;
 wire \u_rf.reg3_q[0] ;
 wire \u_rf.reg3_q[10] ;
 wire \u_rf.reg3_q[11] ;
 wire \u_rf.reg3_q[12] ;
 wire \u_rf.reg3_q[13] ;
 wire \u_rf.reg3_q[14] ;
 wire \u_rf.reg3_q[15] ;
 wire \u_rf.reg3_q[16] ;
 wire \u_rf.reg3_q[17] ;
 wire \u_rf.reg3_q[18] ;
 wire \u_rf.reg3_q[19] ;
 wire \u_rf.reg3_q[1] ;
 wire \u_rf.reg3_q[20] ;
 wire \u_rf.reg3_q[21] ;
 wire \u_rf.reg3_q[22] ;
 wire \u_rf.reg3_q[23] ;
 wire \u_rf.reg3_q[24] ;
 wire \u_rf.reg3_q[25] ;
 wire \u_rf.reg3_q[26] ;
 wire \u_rf.reg3_q[27] ;
 wire \u_rf.reg3_q[28] ;
 wire \u_rf.reg3_q[29] ;
 wire \u_rf.reg3_q[2] ;
 wire \u_rf.reg3_q[30] ;
 wire \u_rf.reg3_q[31] ;
 wire \u_rf.reg3_q[3] ;
 wire \u_rf.reg3_q[4] ;
 wire \u_rf.reg3_q[5] ;
 wire \u_rf.reg3_q[6] ;
 wire \u_rf.reg3_q[7] ;
 wire \u_rf.reg3_q[8] ;
 wire \u_rf.reg3_q[9] ;
 wire \u_rf.reg4_q[0] ;
 wire \u_rf.reg4_q[10] ;
 wire \u_rf.reg4_q[11] ;
 wire \u_rf.reg4_q[12] ;
 wire \u_rf.reg4_q[13] ;
 wire \u_rf.reg4_q[14] ;
 wire \u_rf.reg4_q[15] ;
 wire \u_rf.reg4_q[16] ;
 wire \u_rf.reg4_q[17] ;
 wire \u_rf.reg4_q[18] ;
 wire \u_rf.reg4_q[19] ;
 wire \u_rf.reg4_q[1] ;
 wire \u_rf.reg4_q[20] ;
 wire \u_rf.reg4_q[21] ;
 wire \u_rf.reg4_q[22] ;
 wire \u_rf.reg4_q[23] ;
 wire \u_rf.reg4_q[24] ;
 wire \u_rf.reg4_q[25] ;
 wire \u_rf.reg4_q[26] ;
 wire \u_rf.reg4_q[27] ;
 wire \u_rf.reg4_q[28] ;
 wire \u_rf.reg4_q[29] ;
 wire \u_rf.reg4_q[2] ;
 wire \u_rf.reg4_q[30] ;
 wire \u_rf.reg4_q[31] ;
 wire \u_rf.reg4_q[3] ;
 wire \u_rf.reg4_q[4] ;
 wire \u_rf.reg4_q[5] ;
 wire \u_rf.reg4_q[6] ;
 wire \u_rf.reg4_q[7] ;
 wire \u_rf.reg4_q[8] ;
 wire \u_rf.reg4_q[9] ;
 wire \u_rf.reg5_q[0] ;
 wire \u_rf.reg5_q[10] ;
 wire \u_rf.reg5_q[11] ;
 wire \u_rf.reg5_q[12] ;
 wire \u_rf.reg5_q[13] ;
 wire \u_rf.reg5_q[14] ;
 wire \u_rf.reg5_q[15] ;
 wire \u_rf.reg5_q[16] ;
 wire \u_rf.reg5_q[17] ;
 wire \u_rf.reg5_q[18] ;
 wire \u_rf.reg5_q[19] ;
 wire \u_rf.reg5_q[1] ;
 wire \u_rf.reg5_q[20] ;
 wire \u_rf.reg5_q[21] ;
 wire \u_rf.reg5_q[22] ;
 wire \u_rf.reg5_q[23] ;
 wire \u_rf.reg5_q[24] ;
 wire \u_rf.reg5_q[25] ;
 wire \u_rf.reg5_q[26] ;
 wire \u_rf.reg5_q[27] ;
 wire \u_rf.reg5_q[28] ;
 wire \u_rf.reg5_q[29] ;
 wire \u_rf.reg5_q[2] ;
 wire \u_rf.reg5_q[30] ;
 wire \u_rf.reg5_q[31] ;
 wire \u_rf.reg5_q[3] ;
 wire \u_rf.reg5_q[4] ;
 wire \u_rf.reg5_q[5] ;
 wire \u_rf.reg5_q[6] ;
 wire \u_rf.reg5_q[7] ;
 wire \u_rf.reg5_q[8] ;
 wire \u_rf.reg5_q[9] ;
 wire \u_rf.reg6_q[0] ;
 wire \u_rf.reg6_q[10] ;
 wire \u_rf.reg6_q[11] ;
 wire \u_rf.reg6_q[12] ;
 wire \u_rf.reg6_q[13] ;
 wire \u_rf.reg6_q[14] ;
 wire \u_rf.reg6_q[15] ;
 wire \u_rf.reg6_q[16] ;
 wire \u_rf.reg6_q[17] ;
 wire \u_rf.reg6_q[18] ;
 wire \u_rf.reg6_q[19] ;
 wire \u_rf.reg6_q[1] ;
 wire \u_rf.reg6_q[20] ;
 wire \u_rf.reg6_q[21] ;
 wire \u_rf.reg6_q[22] ;
 wire \u_rf.reg6_q[23] ;
 wire \u_rf.reg6_q[24] ;
 wire \u_rf.reg6_q[25] ;
 wire \u_rf.reg6_q[26] ;
 wire \u_rf.reg6_q[27] ;
 wire \u_rf.reg6_q[28] ;
 wire \u_rf.reg6_q[29] ;
 wire \u_rf.reg6_q[2] ;
 wire \u_rf.reg6_q[30] ;
 wire \u_rf.reg6_q[31] ;
 wire \u_rf.reg6_q[3] ;
 wire \u_rf.reg6_q[4] ;
 wire \u_rf.reg6_q[5] ;
 wire \u_rf.reg6_q[6] ;
 wire \u_rf.reg6_q[7] ;
 wire \u_rf.reg6_q[8] ;
 wire \u_rf.reg6_q[9] ;
 wire \u_rf.reg7_q[0] ;
 wire \u_rf.reg7_q[10] ;
 wire \u_rf.reg7_q[11] ;
 wire \u_rf.reg7_q[12] ;
 wire \u_rf.reg7_q[13] ;
 wire \u_rf.reg7_q[14] ;
 wire \u_rf.reg7_q[15] ;
 wire \u_rf.reg7_q[16] ;
 wire \u_rf.reg7_q[17] ;
 wire \u_rf.reg7_q[18] ;
 wire \u_rf.reg7_q[19] ;
 wire \u_rf.reg7_q[1] ;
 wire \u_rf.reg7_q[20] ;
 wire \u_rf.reg7_q[21] ;
 wire \u_rf.reg7_q[22] ;
 wire \u_rf.reg7_q[23] ;
 wire \u_rf.reg7_q[24] ;
 wire \u_rf.reg7_q[25] ;
 wire \u_rf.reg7_q[26] ;
 wire \u_rf.reg7_q[27] ;
 wire \u_rf.reg7_q[28] ;
 wire \u_rf.reg7_q[29] ;
 wire \u_rf.reg7_q[2] ;
 wire \u_rf.reg7_q[30] ;
 wire \u_rf.reg7_q[31] ;
 wire \u_rf.reg7_q[3] ;
 wire \u_rf.reg7_q[4] ;
 wire \u_rf.reg7_q[5] ;
 wire \u_rf.reg7_q[6] ;
 wire \u_rf.reg7_q[7] ;
 wire \u_rf.reg7_q[8] ;
 wire \u_rf.reg7_q[9] ;
 wire \u_rf.reg8_q[0] ;
 wire \u_rf.reg8_q[10] ;
 wire \u_rf.reg8_q[11] ;
 wire \u_rf.reg8_q[12] ;
 wire \u_rf.reg8_q[13] ;
 wire \u_rf.reg8_q[14] ;
 wire \u_rf.reg8_q[15] ;
 wire \u_rf.reg8_q[16] ;
 wire \u_rf.reg8_q[17] ;
 wire \u_rf.reg8_q[18] ;
 wire \u_rf.reg8_q[19] ;
 wire \u_rf.reg8_q[1] ;
 wire \u_rf.reg8_q[20] ;
 wire \u_rf.reg8_q[21] ;
 wire \u_rf.reg8_q[22] ;
 wire \u_rf.reg8_q[23] ;
 wire \u_rf.reg8_q[24] ;
 wire \u_rf.reg8_q[25] ;
 wire \u_rf.reg8_q[26] ;
 wire \u_rf.reg8_q[27] ;
 wire \u_rf.reg8_q[28] ;
 wire \u_rf.reg8_q[29] ;
 wire \u_rf.reg8_q[2] ;
 wire \u_rf.reg8_q[30] ;
 wire \u_rf.reg8_q[31] ;
 wire \u_rf.reg8_q[3] ;
 wire \u_rf.reg8_q[4] ;
 wire \u_rf.reg8_q[5] ;
 wire \u_rf.reg8_q[6] ;
 wire \u_rf.reg8_q[7] ;
 wire \u_rf.reg8_q[8] ;
 wire \u_rf.reg8_q[9] ;
 wire \u_rf.reg9_q[0] ;
 wire \u_rf.reg9_q[10] ;
 wire \u_rf.reg9_q[11] ;
 wire \u_rf.reg9_q[12] ;
 wire \u_rf.reg9_q[13] ;
 wire \u_rf.reg9_q[14] ;
 wire \u_rf.reg9_q[15] ;
 wire \u_rf.reg9_q[16] ;
 wire \u_rf.reg9_q[17] ;
 wire \u_rf.reg9_q[18] ;
 wire \u_rf.reg9_q[19] ;
 wire \u_rf.reg9_q[1] ;
 wire \u_rf.reg9_q[20] ;
 wire \u_rf.reg9_q[21] ;
 wire \u_rf.reg9_q[22] ;
 wire \u_rf.reg9_q[23] ;
 wire \u_rf.reg9_q[24] ;
 wire \u_rf.reg9_q[25] ;
 wire \u_rf.reg9_q[26] ;
 wire \u_rf.reg9_q[27] ;
 wire \u_rf.reg9_q[28] ;
 wire \u_rf.reg9_q[29] ;
 wire \u_rf.reg9_q[2] ;
 wire \u_rf.reg9_q[30] ;
 wire \u_rf.reg9_q[31] ;
 wire \u_rf.reg9_q[3] ;
 wire \u_rf.reg9_q[4] ;
 wire \u_rf.reg9_q[5] ;
 wire \u_rf.reg9_q[6] ;
 wire \u_rf.reg9_q[7] ;
 wire \u_rf.reg9_q[8] ;
 wire \u_rf.reg9_q[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;

 sky130_fd_sc_hd__nor2_4 _05729_ (.A(\u_exe.flush_v_dly1_q ),
    .B(\u_decod.flush_v ),
    .Y(_01056_));
 sky130_fd_sc_hd__nand2_2 _05730_ (.A(\u_decod.instr_unit_q[3] ),
    .B(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__inv_2 _05731_ (.A(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__buf_2 _05732_ (.A(_01058_),
    .X(_01059_));
 sky130_fd_sc_hd__buf_4 _05733_ (.A(_01059_),
    .X(net133));
 sky130_fd_sc_hd__xor2_2 _05734_ (.A(\u_decod.branch_imm_q_o[1] ),
    .B(\u_decod.rs1_data_q[1] ),
    .X(_01060_));
 sky130_fd_sc_hd__clkbuf_4 _05735_ (.A(\u_decod.rs1_data_q[0] ),
    .X(_01061_));
 sky130_fd_sc_hd__nand2_1 _05736_ (.A(\u_decod.branch_imm_q_o[0] ),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__xnor2_2 _05737_ (.A(_01060_),
    .B(_01062_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand2_1 _05738_ (.A(_01058_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__inv_2 _05739_ (.A(_01064_),
    .Y(net112));
 sky130_fd_sc_hd__or2_1 _05740_ (.A(\u_decod.branch_imm_q_o[0] ),
    .B(_01061_),
    .X(_01065_));
 sky130_fd_sc_hd__nand2_1 _05741_ (.A(_01062_),
    .B(_01065_),
    .Y(_01066_));
 sky130_fd_sc_hd__or2_1 _05742_ (.A(_01057_),
    .B(_01066_),
    .X(_01067_));
 sky130_fd_sc_hd__inv_2 _05743_ (.A(_01067_),
    .Y(net101));
 sky130_fd_sc_hd__nand3b_1 _05744_ (.A_N(\u_decod.dec0.instr_i[4] ),
    .B(\u_decod.dec0.instr_i[5] ),
    .C(\u_decod.dec0.instr_i[6] ),
    .Y(_01068_));
 sky130_fd_sc_hd__nand3_1 _05745_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(\u_decod.dec0.instr_i[1] ),
    .C(\u_decod.dec0.instr_i[2] ),
    .Y(_01069_));
 sky130_fd_sc_hd__or2_1 _05746_ (.A(_01068_),
    .B(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__nor2_1 _05747_ (.A(\u_decod.dec0.instr_i[3] ),
    .B(_01070_),
    .Y(\u_decod.dec0.jalr ));
 sky130_fd_sc_hd__clkbuf_2 _05748_ (.A(\u_decod.dec0.funct3[0] ),
    .X(_01071_));
 sky130_fd_sc_hd__inv_2 _05749_ (.A(\u_decod.dec0.instr_i[3] ),
    .Y(_01072_));
 sky130_fd_sc_hd__and3b_1 _05750_ (.A_N(\u_decod.dec0.instr_i[2] ),
    .B(\u_decod.dec0.instr_i[1] ),
    .C(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__clkbuf_2 _05751_ (.A(_01073_),
    .X(_01074_));
 sky130_fd_sc_hd__and3_2 _05752_ (.A(\u_decod.dec0.instr_i[4] ),
    .B(\u_decod.dec0.instr_i[5] ),
    .C(_01074_),
    .X(_01075_));
 sky130_fd_sc_hd__inv_2 _05753_ (.A(\u_decod.dec0.funct3[1] ),
    .Y(_01076_));
 sky130_fd_sc_hd__nand2b_1 _05754_ (.A_N(\u_decod.dec0.funct3[2] ),
    .B(\u_decod.dec0.instr_i[0] ),
    .Y(_01077_));
 sky130_fd_sc_hd__nor2_1 _05755_ (.A(_01076_),
    .B(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__buf_4 _05756_ (.A(\u_decod.dec0.funct7[5] ),
    .X(_01079_));
 sky130_fd_sc_hd__clkbuf_2 _05757_ (.A(\u_decod.dec0.instr_i[6] ),
    .X(_01080_));
 sky130_fd_sc_hd__or2_1 _05758_ (.A(\u_decod.dec0.funct7[1] ),
    .B(\u_decod.dec0.funct7[0] ),
    .X(_01081_));
 sky130_fd_sc_hd__or4_1 _05759_ (.A(\u_decod.dec0.funct7[3] ),
    .B(\u_decod.dec0.funct7[2] ),
    .C(\u_decod.dec0.funct7[4] ),
    .D(_01081_),
    .X(_01082_));
 sky130_fd_sc_hd__or3_1 _05760_ (.A(_01080_),
    .B(\u_decod.dec0.funct7[6] ),
    .C(_01082_),
    .X(_01083_));
 sky130_fd_sc_hd__nor2_1 _05761_ (.A(_01079_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__or2_1 _05762_ (.A(_01076_),
    .B(_01077_),
    .X(_01085_));
 sky130_fd_sc_hd__and2_1 _05763_ (.A(\u_decod.dec0.instr_i[4] ),
    .B(_01074_),
    .X(_01086_));
 sky130_fd_sc_hd__nor2_1 _05764_ (.A(\u_decod.dec0.instr_i[6] ),
    .B(\u_decod.dec0.instr_i[5] ),
    .Y(_01087_));
 sky130_fd_sc_hd__nand2_1 _05765_ (.A(_01086_),
    .B(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__nor2_1 _05766_ (.A(_01085_),
    .B(_01088_),
    .Y(_01089_));
 sky130_fd_sc_hd__and2b_2 _05767_ (.A_N(_01068_),
    .B(_01074_),
    .X(_01090_));
 sky130_fd_sc_hd__and3_1 _05768_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(\u_decod.dec0.funct3[1] ),
    .C(\u_decod.dec0.funct3[2] ),
    .X(_01091_));
 sky130_fd_sc_hd__and2b_1 _05769_ (.A_N(\u_decod.dec0.instr_i[4] ),
    .B(_01087_),
    .X(_01092_));
 sky130_fd_sc_hd__and2_1 _05770_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(\u_decod.dec0.funct3[2] ),
    .X(_01093_));
 sky130_fd_sc_hd__and2_1 _05771_ (.A(_01076_),
    .B(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__and3_1 _05772_ (.A(_01074_),
    .B(_01092_),
    .C(_01094_),
    .X(_01095_));
 sky130_fd_sc_hd__a221o_1 _05773_ (.A1(_01071_),
    .A2(_01089_),
    .B1(_01090_),
    .B2(_01091_),
    .C1(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__a41o_1 _05774_ (.A1(_01071_),
    .A2(_01075_),
    .A3(_01078_),
    .A4(_01084_),
    .B1(_01096_),
    .X(_01097_));
 sky130_fd_sc_hd__clkbuf_2 _05775_ (.A(_01097_),
    .X(\u_decod.dec0.unsign_extension ));
 sky130_fd_sc_hd__and2b_1 _05776_ (.A_N(\u_decod.flush_v ),
    .B(net361),
    .X(_01098_));
 sky130_fd_sc_hd__buf_4 _05777_ (.A(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__nor2b_2 _05778_ (.A(\u_ifetch.reset_n_q ),
    .B_N(net369),
    .Y(_01100_));
 sky130_fd_sc_hd__buf_2 _05779_ (.A(_01100_),
    .X(_01101_));
 sky130_fd_sc_hd__and3_1 _05780_ (.A(\u_decod.flush_v ),
    .B(net360),
    .C(\u_exe.pc_data_q[0] ),
    .X(_01102_));
 sky130_fd_sc_hd__a221o_1 _05781_ (.A1(\u_decod.pc0_q_i[0] ),
    .A2(_01099_),
    .B1(_01101_),
    .B2(net65),
    .C1(_01102_),
    .X(net134));
 sky130_fd_sc_hd__and3_1 _05782_ (.A(\u_decod.flush_v ),
    .B(net360),
    .C(\u_exe.pc_data_q[1] ),
    .X(_01103_));
 sky130_fd_sc_hd__a221o_1 _05783_ (.A1(\u_decod.pc0_q_i[1] ),
    .A2(_01099_),
    .B1(_01101_),
    .B2(net76),
    .C1(_01103_),
    .X(net145));
 sky130_fd_sc_hd__and2_1 _05784_ (.A(\u_decod.flush_v ),
    .B(net361),
    .X(_01104_));
 sky130_fd_sc_hd__clkbuf_4 _05785_ (.A(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__buf_2 _05786_ (.A(_01098_),
    .X(_01106_));
 sky130_fd_sc_hd__and2b_1 _05787_ (.A_N(\u_decod.pc0_q_i[2] ),
    .B(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__a221o_1 _05788_ (.A1(\u_exe.pc_data_q[2] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net87),
    .C1(_01107_),
    .X(net156));
 sky130_fd_sc_hd__a21boi_1 _05789_ (.A1(\u_decod.pc0_q_i[2] ),
    .A2(\u_decod.pc0_q_i[3] ),
    .B1_N(_01098_),
    .Y(_01108_));
 sky130_fd_sc_hd__o21a_1 _05790_ (.A1(\u_decod.pc0_q_i[2] ),
    .A2(\u_decod.pc0_q_i[3] ),
    .B1(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__a221o_2 _05791_ (.A1(\u_exe.pc_data_q[3] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net90),
    .C1(_01109_),
    .X(net159));
 sky130_fd_sc_hd__and3_1 _05792_ (.A(\u_decod.pc0_q_i[2] ),
    .B(\u_decod.pc0_q_i[3] ),
    .C(\u_decod.pc0_q_i[4] ),
    .X(_01110_));
 sky130_fd_sc_hd__a21o_1 _05793_ (.A1(\u_decod.pc0_q_i[2] ),
    .A2(\u_decod.pc0_q_i[3] ),
    .B1(\u_decod.pc0_q_i[4] ),
    .X(_01111_));
 sky130_fd_sc_hd__and3b_1 _05794_ (.A_N(_01110_),
    .B(_01106_),
    .C(_01111_),
    .X(_01112_));
 sky130_fd_sc_hd__a221o_2 _05795_ (.A1(\u_exe.pc_data_q[4] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net91),
    .C1(_01112_),
    .X(net160));
 sky130_fd_sc_hd__and4_1 _05796_ (.A(\u_decod.pc0_q_i[2] ),
    .B(\u_decod.pc0_q_i[3] ),
    .C(\u_decod.pc0_q_i[4] ),
    .D(\u_decod.pc0_q_i[5] ),
    .X(_01113_));
 sky130_fd_sc_hd__or2_1 _05797_ (.A(\u_decod.pc0_q_i[5] ),
    .B(_01110_),
    .X(_01114_));
 sky130_fd_sc_hd__and3b_1 _05798_ (.A_N(_01113_),
    .B(_01106_),
    .C(_01114_),
    .X(_01115_));
 sky130_fd_sc_hd__a221o_1 _05799_ (.A1(\u_exe.pc_data_q[5] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net92),
    .C1(_01115_),
    .X(net161));
 sky130_fd_sc_hd__or2_1 _05800_ (.A(\u_decod.pc0_q_i[6] ),
    .B(_01113_),
    .X(_01116_));
 sky130_fd_sc_hd__nand2_1 _05801_ (.A(\u_decod.pc0_q_i[6] ),
    .B(_01113_),
    .Y(_01117_));
 sky130_fd_sc_hd__clkbuf_4 _05802_ (.A(_01104_),
    .X(_01118_));
 sky130_fd_sc_hd__clkbuf_4 _05803_ (.A(_01100_),
    .X(_01119_));
 sky130_fd_sc_hd__a22o_1 _05804_ (.A1(\u_exe.pc_data_q[6] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net93),
    .X(_01120_));
 sky130_fd_sc_hd__a31o_2 _05805_ (.A1(_01099_),
    .A2(_01116_),
    .A3(_01117_),
    .B1(_01120_),
    .X(net162));
 sky130_fd_sc_hd__and3_1 _05806_ (.A(\u_decod.pc0_q_i[6] ),
    .B(\u_decod.pc0_q_i[7] ),
    .C(_01113_),
    .X(_01121_));
 sky130_fd_sc_hd__a21o_1 _05807_ (.A1(\u_decod.pc0_q_i[6] ),
    .A2(_01113_),
    .B1(\u_decod.pc0_q_i[7] ),
    .X(_01122_));
 sky130_fd_sc_hd__and3b_1 _05808_ (.A_N(_01121_),
    .B(_01106_),
    .C(_01122_),
    .X(_01123_));
 sky130_fd_sc_hd__a221o_1 _05809_ (.A1(\u_exe.pc_data_q[7] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net94),
    .C1(_01123_),
    .X(net163));
 sky130_fd_sc_hd__and4_1 _05810_ (.A(\u_decod.pc0_q_i[6] ),
    .B(\u_decod.pc0_q_i[7] ),
    .C(\u_decod.pc0_q_i[8] ),
    .D(_01113_),
    .X(_01124_));
 sky130_fd_sc_hd__or2_1 _05811_ (.A(\u_decod.pc0_q_i[8] ),
    .B(_01121_),
    .X(_01125_));
 sky130_fd_sc_hd__and3b_1 _05812_ (.A_N(_01124_),
    .B(_01106_),
    .C(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__a221o_1 _05813_ (.A1(\u_exe.pc_data_q[8] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net95),
    .C1(_01126_),
    .X(net164));
 sky130_fd_sc_hd__o21ai_1 _05814_ (.A1(\u_decod.pc0_q_i[9] ),
    .A2(_01124_),
    .B1(_01106_),
    .Y(_01127_));
 sky130_fd_sc_hd__a21oi_1 _05815_ (.A1(\u_decod.pc0_q_i[9] ),
    .A2(_01124_),
    .B1(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__a221o_1 _05816_ (.A1(\u_exe.pc_data_q[9] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net96),
    .C1(_01128_),
    .X(net165));
 sky130_fd_sc_hd__and3_1 _05817_ (.A(\u_decod.pc0_q_i[9] ),
    .B(\u_decod.pc0_q_i[10] ),
    .C(_01124_),
    .X(_01129_));
 sky130_fd_sc_hd__a21o_1 _05818_ (.A1(\u_decod.pc0_q_i[9] ),
    .A2(_01124_),
    .B1(\u_decod.pc0_q_i[10] ),
    .X(_01130_));
 sky130_fd_sc_hd__and3b_1 _05819_ (.A_N(_01129_),
    .B(_01106_),
    .C(_01130_),
    .X(_01131_));
 sky130_fd_sc_hd__a221o_1 _05820_ (.A1(\u_exe.pc_data_q[10] ),
    .A2(_01105_),
    .B1(_01101_),
    .B2(net66),
    .C1(_01131_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 _05821_ (.A(_01100_),
    .X(_01132_));
 sky130_fd_sc_hd__and2_1 _05822_ (.A(\u_decod.pc0_q_i[11] ),
    .B(_01129_),
    .X(_01133_));
 sky130_fd_sc_hd__or2_1 _05823_ (.A(\u_decod.pc0_q_i[11] ),
    .B(_01129_),
    .X(_01134_));
 sky130_fd_sc_hd__and3b_1 _05824_ (.A_N(_01133_),
    .B(_01106_),
    .C(_01134_),
    .X(_01135_));
 sky130_fd_sc_hd__a221o_1 _05825_ (.A1(\u_exe.pc_data_q[11] ),
    .A2(_01105_),
    .B1(_01132_),
    .B2(net67),
    .C1(_01135_),
    .X(net136));
 sky130_fd_sc_hd__or2_1 _05826_ (.A(\u_decod.pc0_q_i[12] ),
    .B(_01133_),
    .X(_01136_));
 sky130_fd_sc_hd__nand2_1 _05827_ (.A(\u_decod.pc0_q_i[12] ),
    .B(_01133_),
    .Y(_01137_));
 sky130_fd_sc_hd__a22o_1 _05828_ (.A1(\u_exe.pc_data_q[12] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net68),
    .X(_01138_));
 sky130_fd_sc_hd__a31o_1 _05829_ (.A1(_01099_),
    .A2(_01136_),
    .A3(_01137_),
    .B1(_01138_),
    .X(net137));
 sky130_fd_sc_hd__and3_1 _05830_ (.A(\u_decod.pc0_q_i[12] ),
    .B(\u_decod.pc0_q_i[13] ),
    .C(_01133_),
    .X(_01139_));
 sky130_fd_sc_hd__a31o_1 _05831_ (.A1(\u_decod.pc0_q_i[11] ),
    .A2(\u_decod.pc0_q_i[12] ),
    .A3(_01129_),
    .B1(\u_decod.pc0_q_i[13] ),
    .X(_01140_));
 sky130_fd_sc_hd__and3b_1 _05832_ (.A_N(_01139_),
    .B(_01106_),
    .C(_01140_),
    .X(_01141_));
 sky130_fd_sc_hd__a221o_1 _05833_ (.A1(\u_exe.pc_data_q[13] ),
    .A2(_01105_),
    .B1(_01132_),
    .B2(net69),
    .C1(_01141_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 _05834_ (.A(_01104_),
    .X(_01142_));
 sky130_fd_sc_hd__and2_1 _05835_ (.A(\u_decod.pc0_q_i[14] ),
    .B(_01139_),
    .X(_01143_));
 sky130_fd_sc_hd__buf_2 _05836_ (.A(_01098_),
    .X(_01144_));
 sky130_fd_sc_hd__or2_1 _05837_ (.A(\u_decod.pc0_q_i[14] ),
    .B(_01139_),
    .X(_01145_));
 sky130_fd_sc_hd__and3b_1 _05838_ (.A_N(_01143_),
    .B(_01144_),
    .C(_01145_),
    .X(_01146_));
 sky130_fd_sc_hd__a221o_1 _05839_ (.A1(\u_exe.pc_data_q[14] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net70),
    .C1(_01146_),
    .X(net139));
 sky130_fd_sc_hd__or2_1 _05840_ (.A(\u_decod.pc0_q_i[15] ),
    .B(_01143_),
    .X(_01147_));
 sky130_fd_sc_hd__nand2_1 _05841_ (.A(\u_decod.pc0_q_i[15] ),
    .B(_01143_),
    .Y(_01148_));
 sky130_fd_sc_hd__a22o_1 _05842_ (.A1(\u_exe.pc_data_q[15] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net71),
    .X(_01149_));
 sky130_fd_sc_hd__a31o_1 _05843_ (.A1(_01099_),
    .A2(_01147_),
    .A3(_01148_),
    .B1(_01149_),
    .X(net140));
 sky130_fd_sc_hd__and3_1 _05844_ (.A(\u_decod.pc0_q_i[15] ),
    .B(\u_decod.pc0_q_i[16] ),
    .C(_01143_),
    .X(_01150_));
 sky130_fd_sc_hd__a31o_1 _05845_ (.A1(\u_decod.pc0_q_i[14] ),
    .A2(\u_decod.pc0_q_i[15] ),
    .A3(_01139_),
    .B1(\u_decod.pc0_q_i[16] ),
    .X(_01151_));
 sky130_fd_sc_hd__and3b_1 _05846_ (.A_N(_01150_),
    .B(_01144_),
    .C(_01151_),
    .X(_01152_));
 sky130_fd_sc_hd__a221o_1 _05847_ (.A1(\u_exe.pc_data_q[16] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net72),
    .C1(_01152_),
    .X(net141));
 sky130_fd_sc_hd__and2_1 _05848_ (.A(\u_decod.pc0_q_i[17] ),
    .B(_01150_),
    .X(_01153_));
 sky130_fd_sc_hd__or2_1 _05849_ (.A(\u_decod.pc0_q_i[17] ),
    .B(_01150_),
    .X(_01154_));
 sky130_fd_sc_hd__and3b_1 _05850_ (.A_N(_01153_),
    .B(_01144_),
    .C(_01154_),
    .X(_01155_));
 sky130_fd_sc_hd__a221o_1 _05851_ (.A1(\u_exe.pc_data_q[17] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net73),
    .C1(_01155_),
    .X(net142));
 sky130_fd_sc_hd__or2_1 _05852_ (.A(\u_decod.pc0_q_i[18] ),
    .B(_01153_),
    .X(_01156_));
 sky130_fd_sc_hd__nand2_1 _05853_ (.A(\u_decod.pc0_q_i[18] ),
    .B(_01153_),
    .Y(_01157_));
 sky130_fd_sc_hd__a22o_1 _05854_ (.A1(\u_exe.pc_data_q[18] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net74),
    .X(_01158_));
 sky130_fd_sc_hd__a31o_1 _05855_ (.A1(_01099_),
    .A2(_01156_),
    .A3(_01157_),
    .B1(_01158_),
    .X(net143));
 sky130_fd_sc_hd__and3_1 _05856_ (.A(\u_decod.pc0_q_i[18] ),
    .B(\u_decod.pc0_q_i[19] ),
    .C(_01153_),
    .X(_01159_));
 sky130_fd_sc_hd__a31o_1 _05857_ (.A1(\u_decod.pc0_q_i[17] ),
    .A2(\u_decod.pc0_q_i[18] ),
    .A3(_01150_),
    .B1(\u_decod.pc0_q_i[19] ),
    .X(_01160_));
 sky130_fd_sc_hd__and3b_1 _05858_ (.A_N(_01159_),
    .B(_01144_),
    .C(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__a221o_1 _05859_ (.A1(\u_exe.pc_data_q[19] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net75),
    .C1(_01161_),
    .X(net144));
 sky130_fd_sc_hd__and2_1 _05860_ (.A(\u_decod.pc0_q_i[20] ),
    .B(_01159_),
    .X(_01162_));
 sky130_fd_sc_hd__or2_1 _05861_ (.A(\u_decod.pc0_q_i[20] ),
    .B(_01159_),
    .X(_01163_));
 sky130_fd_sc_hd__and3b_1 _05862_ (.A_N(_01162_),
    .B(_01144_),
    .C(_01163_),
    .X(_01164_));
 sky130_fd_sc_hd__a221o_1 _05863_ (.A1(\u_exe.pc_data_q[20] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net77),
    .C1(_01164_),
    .X(net146));
 sky130_fd_sc_hd__or2_1 _05864_ (.A(\u_decod.pc0_q_i[21] ),
    .B(_01162_),
    .X(_01165_));
 sky130_fd_sc_hd__nand2_1 _05865_ (.A(\u_decod.pc0_q_i[21] ),
    .B(_01162_),
    .Y(_01166_));
 sky130_fd_sc_hd__a22o_1 _05866_ (.A1(\u_exe.pc_data_q[21] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net78),
    .X(_01167_));
 sky130_fd_sc_hd__a31o_1 _05867_ (.A1(_01099_),
    .A2(_01165_),
    .A3(_01166_),
    .B1(_01167_),
    .X(net147));
 sky130_fd_sc_hd__and3_1 _05868_ (.A(\u_decod.pc0_q_i[21] ),
    .B(\u_decod.pc0_q_i[22] ),
    .C(_01162_),
    .X(_01168_));
 sky130_fd_sc_hd__a31o_1 _05869_ (.A1(\u_decod.pc0_q_i[20] ),
    .A2(\u_decod.pc0_q_i[21] ),
    .A3(_01159_),
    .B1(\u_decod.pc0_q_i[22] ),
    .X(_01169_));
 sky130_fd_sc_hd__and3b_1 _05870_ (.A_N(_01168_),
    .B(_01144_),
    .C(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__a221o_1 _05871_ (.A1(\u_exe.pc_data_q[22] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net79),
    .C1(_01170_),
    .X(net148));
 sky130_fd_sc_hd__and2_1 _05872_ (.A(\u_decod.pc0_q_i[23] ),
    .B(_01168_),
    .X(_01171_));
 sky130_fd_sc_hd__or2_1 _05873_ (.A(\u_decod.pc0_q_i[23] ),
    .B(_01168_),
    .X(_01172_));
 sky130_fd_sc_hd__and3b_1 _05874_ (.A_N(_01171_),
    .B(_01144_),
    .C(_01172_),
    .X(_01173_));
 sky130_fd_sc_hd__a221o_1 _05875_ (.A1(\u_exe.pc_data_q[23] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net80),
    .C1(_01173_),
    .X(net149));
 sky130_fd_sc_hd__or2_1 _05876_ (.A(\u_decod.pc0_q_i[24] ),
    .B(_01171_),
    .X(_01174_));
 sky130_fd_sc_hd__nand2_1 _05877_ (.A(\u_decod.pc0_q_i[24] ),
    .B(_01171_),
    .Y(_01175_));
 sky130_fd_sc_hd__a22o_1 _05878_ (.A1(\u_exe.pc_data_q[24] ),
    .A2(_01118_),
    .B1(_01100_),
    .B2(net81),
    .X(_01176_));
 sky130_fd_sc_hd__a31o_1 _05879_ (.A1(_01099_),
    .A2(_01174_),
    .A3(_01175_),
    .B1(_01176_),
    .X(net150));
 sky130_fd_sc_hd__and3_1 _05880_ (.A(\u_decod.pc0_q_i[24] ),
    .B(\u_decod.pc0_q_i[25] ),
    .C(_01171_),
    .X(_01177_));
 sky130_fd_sc_hd__a31o_1 _05881_ (.A1(\u_decod.pc0_q_i[23] ),
    .A2(\u_decod.pc0_q_i[24] ),
    .A3(_01168_),
    .B1(\u_decod.pc0_q_i[25] ),
    .X(_01178_));
 sky130_fd_sc_hd__and3b_1 _05882_ (.A_N(_01177_),
    .B(_01144_),
    .C(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__a221o_1 _05883_ (.A1(\u_exe.pc_data_q[25] ),
    .A2(_01142_),
    .B1(_01132_),
    .B2(net82),
    .C1(_01179_),
    .X(net151));
 sky130_fd_sc_hd__and2_1 _05884_ (.A(\u_decod.pc0_q_i[26] ),
    .B(_01177_),
    .X(_01180_));
 sky130_fd_sc_hd__or2_1 _05885_ (.A(\u_decod.pc0_q_i[26] ),
    .B(_01177_),
    .X(_01181_));
 sky130_fd_sc_hd__and3b_1 _05886_ (.A_N(_01180_),
    .B(_01144_),
    .C(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__a221o_1 _05887_ (.A1(\u_exe.pc_data_q[26] ),
    .A2(_01142_),
    .B1(_01119_),
    .B2(net83),
    .C1(_01182_),
    .X(net152));
 sky130_fd_sc_hd__or2_1 _05888_ (.A(\u_decod.pc0_q_i[27] ),
    .B(_01180_),
    .X(_01183_));
 sky130_fd_sc_hd__nand2_1 _05889_ (.A(\u_decod.pc0_q_i[27] ),
    .B(_01180_),
    .Y(_01184_));
 sky130_fd_sc_hd__a22o_1 _05890_ (.A1(\u_exe.pc_data_q[27] ),
    .A2(_01118_),
    .B1(_01100_),
    .B2(net84),
    .X(_01185_));
 sky130_fd_sc_hd__a31o_1 _05891_ (.A1(_01099_),
    .A2(_01183_),
    .A3(_01184_),
    .B1(_01185_),
    .X(net153));
 sky130_fd_sc_hd__and3_1 _05892_ (.A(\u_decod.pc0_q_i[27] ),
    .B(\u_decod.pc0_q_i[28] ),
    .C(_01180_),
    .X(_01186_));
 sky130_fd_sc_hd__a31o_1 _05893_ (.A1(\u_decod.pc0_q_i[26] ),
    .A2(\u_decod.pc0_q_i[27] ),
    .A3(_01177_),
    .B1(\u_decod.pc0_q_i[28] ),
    .X(_01187_));
 sky130_fd_sc_hd__and3b_1 _05894_ (.A_N(_01186_),
    .B(_01144_),
    .C(_01187_),
    .X(_01188_));
 sky130_fd_sc_hd__a221o_1 _05895_ (.A1(\u_exe.pc_data_q[28] ),
    .A2(_01142_),
    .B1(_01119_),
    .B2(net85),
    .C1(_01188_),
    .X(net154));
 sky130_fd_sc_hd__and2_1 _05896_ (.A(\u_decod.pc0_q_i[29] ),
    .B(_01186_),
    .X(_01189_));
 sky130_fd_sc_hd__o21ai_1 _05897_ (.A1(\u_decod.pc0_q_i[29] ),
    .A2(_01186_),
    .B1(_01099_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _05898_ (.A(_01189_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__a221o_1 _05899_ (.A1(\u_exe.pc_data_q[29] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net86),
    .C1(_01191_),
    .X(net155));
 sky130_fd_sc_hd__and3_1 _05900_ (.A(\u_decod.pc0_q_i[29] ),
    .B(\u_decod.pc0_q_i[30] ),
    .C(_01186_),
    .X(_01192_));
 sky130_fd_sc_hd__or2_1 _05901_ (.A(\u_decod.pc0_q_i[30] ),
    .B(_01189_),
    .X(_01193_));
 sky130_fd_sc_hd__and3b_1 _05902_ (.A_N(_01192_),
    .B(_01098_),
    .C(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a221o_1 _05903_ (.A1(\u_exe.pc_data_q[30] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net88),
    .C1(_01194_),
    .X(net157));
 sky130_fd_sc_hd__o21ai_1 _05904_ (.A1(\u_decod.pc0_q_i[31] ),
    .A2(_01192_),
    .B1(_01106_),
    .Y(_01195_));
 sky130_fd_sc_hd__a21oi_1 _05905_ (.A1(\u_decod.pc0_q_i[31] ),
    .A2(_01192_),
    .B1(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__a221o_1 _05906_ (.A1(\u_exe.pc_data_q[31] ),
    .A2(_01118_),
    .B1(_01119_),
    .B2(net89),
    .C1(_01196_),
    .X(net158));
 sky130_fd_sc_hd__or2_1 _05907_ (.A(\u_decod.dec0.funct3[1] ),
    .B(_01077_),
    .X(_01197_));
 sky130_fd_sc_hd__nor2_1 _05908_ (.A(_01071_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__and2_1 _05909_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(_01074_),
    .X(_01199_));
 sky130_fd_sc_hd__a41o_1 _05910_ (.A1(\u_decod.dec0.instr_i[1] ),
    .A2(\u_decod.dec0.instr_i[3] ),
    .A3(\u_decod.dec0.instr_i[2] ),
    .A4(_01198_),
    .B1(_01199_),
    .X(_01200_));
 sky130_fd_sc_hd__nand2_1 _05911_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(_01074_),
    .Y(_01201_));
 sky130_fd_sc_hd__or3b_1 _05912_ (.A(_01201_),
    .B(_01080_),
    .C_N(\u_decod.dec0.instr_i[4] ),
    .X(_01202_));
 sky130_fd_sc_hd__inv_2 _05913_ (.A(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__a211o_1 _05914_ (.A1(_01092_),
    .A2(_01200_),
    .B1(_01203_),
    .C1(\u_decod.dec0.jalr ),
    .X(_01204_));
 sky130_fd_sc_hd__nor2_1 _05915_ (.A(_01072_),
    .B(_01070_),
    .Y(_01205_));
 sky130_fd_sc_hd__and4bb_4 _05916_ (.A_N(_01069_),
    .B_N(_01080_),
    .C(_01072_),
    .D(\u_decod.dec0.instr_i[4] ),
    .X(_01206_));
 sky130_fd_sc_hd__or2_1 _05917_ (.A(_01205_),
    .B(_01206_),
    .X(_01207_));
 sky130_fd_sc_hd__clkbuf_4 _05918_ (.A(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__or2_1 _05919_ (.A(_01079_),
    .B(_01082_),
    .X(_01209_));
 sky130_fd_sc_hd__or3_1 _05920_ (.A(\u_decod.dec0.funct3[0] ),
    .B(\u_decod.dec0.funct7[6] ),
    .C(\u_decod.dec0.instr_i[20] ),
    .X(_01210_));
 sky130_fd_sc_hd__or4_1 _05921_ (.A(\u_decod.dec0.funct3[1] ),
    .B(\u_decod.dec0.funct3[2] ),
    .C(_01209_),
    .D(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__nand4_1 _05922_ (.A(\u_decod.dec0.instr_i[0] ),
    .B(_01080_),
    .C(_01075_),
    .D(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__or3b_1 _05923_ (.A(_01204_),
    .B(_01208_),
    .C_N(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__clkbuf_2 _05924_ (.A(_01213_),
    .X(\u_decod.dec0.rd_v ));
 sky130_fd_sc_hd__and2_1 _05925_ (.A(\u_decod.dec0.instr_i[7] ),
    .B(\u_decod.dec0.rd_v ),
    .X(_01214_));
 sky130_fd_sc_hd__clkbuf_1 _05926_ (.A(_01214_),
    .X(\u_decod.dec0.rd_o[0] ));
 sky130_fd_sc_hd__and2_1 _05927_ (.A(\u_decod.dec0.instr_i[8] ),
    .B(\u_decod.dec0.rd_v ),
    .X(_01215_));
 sky130_fd_sc_hd__clkbuf_1 _05928_ (.A(_01215_),
    .X(\u_decod.dec0.rd_o[1] ));
 sky130_fd_sc_hd__and2_1 _05929_ (.A(\u_decod.dec0.instr_i[9] ),
    .B(\u_decod.dec0.rd_v ),
    .X(_01216_));
 sky130_fd_sc_hd__clkbuf_1 _05930_ (.A(_01216_),
    .X(\u_decod.dec0.rd_o[2] ));
 sky130_fd_sc_hd__and2_1 _05931_ (.A(\u_decod.dec0.instr_i[10] ),
    .B(\u_decod.dec0.rd_v ),
    .X(_01217_));
 sky130_fd_sc_hd__clkbuf_1 _05932_ (.A(_01217_),
    .X(\u_decod.dec0.rd_o[3] ));
 sky130_fd_sc_hd__and2_1 _05933_ (.A(\u_decod.dec0.instr_i[11] ),
    .B(\u_decod.dec0.rd_v ),
    .X(_01218_));
 sky130_fd_sc_hd__clkbuf_1 _05934_ (.A(_01218_),
    .X(\u_decod.dec0.rd_o[4] ));
 sky130_fd_sc_hd__o21ai_1 _05935_ (.A1(_01068_),
    .A2(_01201_),
    .B1(_01070_),
    .Y(\u_decod.dec0.is_branch ));
 sky130_fd_sc_hd__nor3_1 _05936_ (.A(_01080_),
    .B(\u_decod.dec0.funct7[6] ),
    .C(_01082_),
    .Y(_01219_));
 sky130_fd_sc_hd__and4_1 _05937_ (.A(_01071_),
    .B(_01086_),
    .C(_01219_),
    .D(_01094_),
    .X(_01220_));
 sky130_fd_sc_hd__nor2_1 _05938_ (.A(\u_decod.dec0.funct3[1] ),
    .B(_01077_),
    .Y(_01221_));
 sky130_fd_sc_hd__and4_1 _05939_ (.A(_01071_),
    .B(_01086_),
    .C(_01084_),
    .D(_01221_),
    .X(_01222_));
 sky130_fd_sc_hd__or2_1 _05940_ (.A(_01220_),
    .B(_01222_),
    .X(_01223_));
 sky130_fd_sc_hd__clkbuf_1 _05941_ (.A(_01223_),
    .X(\u_decod.dec0.is_shift ));
 sky130_fd_sc_hd__clkbuf_4 _05942_ (.A(_01206_),
    .X(_01224_));
 sky130_fd_sc_hd__o21bai_1 _05943_ (.A1(_01202_),
    .A2(\u_decod.dec0.is_shift ),
    .B1_N(_01224_),
    .Y(\u_decod.dec0.is_arithm ));
 sky130_fd_sc_hd__nand2_2 _05944_ (.A(\u_decod.dec0.instr_i[5] ),
    .B(_01199_),
    .Y(_01225_));
 sky130_fd_sc_hd__nor2_4 _05945_ (.A(\u_decod.dec0.instr_i[4] ),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__and2b_1 _05946_ (.A_N(_01080_),
    .B(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__a21oi_1 _05947_ (.A1(_01071_),
    .A2(\u_decod.dec0.funct3[1] ),
    .B1(_01077_),
    .Y(_01228_));
 sky130_fd_sc_hd__o211a_1 _05948_ (.A1(_01094_),
    .A2(_01228_),
    .B1(_01074_),
    .C1(_01092_),
    .X(_01229_));
 sky130_fd_sc_hd__or2_1 _05949_ (.A(_01227_),
    .B(_01229_),
    .X(_01230_));
 sky130_fd_sc_hd__clkbuf_1 _05950_ (.A(_01230_),
    .X(\u_decod.dec0.unit_o[3] ));
 sky130_fd_sc_hd__nand2_1 _05951_ (.A(\u_decod.dec0.instr_i[5] ),
    .B(_01086_),
    .Y(_01231_));
 sky130_fd_sc_hd__or3_1 _05952_ (.A(_01080_),
    .B(\u_decod.dec0.funct3[0] ),
    .C(\u_decod.dec0.funct7[6] ),
    .X(_01232_));
 sky130_fd_sc_hd__or4_1 _05953_ (.A(_01231_),
    .B(_01085_),
    .C(_01209_),
    .D(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__inv_2 _05954_ (.A(\u_decod.dec0.funct3[0] ),
    .Y(_01234_));
 sky130_fd_sc_hd__or3_1 _05955_ (.A(_01080_),
    .B(_01234_),
    .C(\u_decod.dec0.funct7[6] ),
    .X(_01235_));
 sky130_fd_sc_hd__or4_1 _05956_ (.A(_01231_),
    .B(_01085_),
    .C(_01209_),
    .D(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__nand3b_2 _05957_ (.A_N(_01089_),
    .B(_01233_),
    .C(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__or2_1 _05958_ (.A(_01205_),
    .B(_01237_),
    .X(_01238_));
 sky130_fd_sc_hd__clkbuf_1 _05959_ (.A(_01238_),
    .X(\u_decod.dec0.operation_o[4] ));
 sky130_fd_sc_hd__inv_2 _05960_ (.A(_01088_),
    .Y(_01239_));
 sky130_fd_sc_hd__a21o_1 _05961_ (.A1(_01075_),
    .A2(_01084_),
    .B1(_01239_),
    .X(_01240_));
 sky130_fd_sc_hd__nor2_1 _05962_ (.A(_01068_),
    .B(_01201_),
    .Y(_01241_));
 sky130_fd_sc_hd__and3_1 _05963_ (.A(_01071_),
    .B(\u_decod.dec0.funct3[2] ),
    .C(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__a31o_1 _05964_ (.A1(_01234_),
    .A2(_01094_),
    .A3(_01240_),
    .B1(_01242_),
    .X(\u_decod.dec0.operation_o[3] ));
 sky130_fd_sc_hd__and2_2 _05965_ (.A(\u_decod.dec0.funct3[2] ),
    .B(_01241_),
    .X(_01243_));
 sky130_fd_sc_hd__and3_1 _05966_ (.A(_01086_),
    .B(_01087_),
    .C(_01091_),
    .X(_01244_));
 sky130_fd_sc_hd__a311o_1 _05967_ (.A1(_01075_),
    .A2(_01084_),
    .A3(_01091_),
    .B1(_01243_),
    .C1(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__a22o_1 _05968_ (.A1(_01079_),
    .A2(_01220_),
    .B1(_01245_),
    .B2(_01234_),
    .X(\u_decod.dec0.operation_o[2] ));
 sky130_fd_sc_hd__o211a_1 _05969_ (.A1(\u_decod.dec0.instr_i[5] ),
    .A2(_01076_),
    .B1(_01086_),
    .C1(_01093_),
    .X(_01246_));
 sky130_fd_sc_hd__a221o_1 _05970_ (.A1(_01090_),
    .A2(_01221_),
    .B1(_01246_),
    .B2(_01084_),
    .C1(_01244_),
    .X(_01247_));
 sky130_fd_sc_hd__a21o_1 _05971_ (.A1(_01071_),
    .A2(_01247_),
    .B1(_01229_),
    .X(\u_decod.dec0.operation_o[1] ));
 sky130_fd_sc_hd__or2_1 _05972_ (.A(_01224_),
    .B(_01222_),
    .X(_01248_));
 sky130_fd_sc_hd__o21a_1 _05973_ (.A1(_01239_),
    .A2(_01090_),
    .B1(_01198_),
    .X(_01249_));
 sky130_fd_sc_hd__and3_1 _05974_ (.A(_01075_),
    .B(_01219_),
    .C(_01198_),
    .X(_01250_));
 sky130_fd_sc_hd__or4_1 _05975_ (.A(_01227_),
    .B(_01248_),
    .C(_01249_),
    .D(_01250_),
    .X(_01251_));
 sky130_fd_sc_hd__clkbuf_1 _05976_ (.A(_01251_),
    .X(\u_decod.dec0.operation_o[0] ));
 sky130_fd_sc_hd__nor2_1 _05977_ (.A(_01080_),
    .B(\u_decod.dec0.instr_i[4] ),
    .Y(_01252_));
 sky130_fd_sc_hd__a31o_1 _05978_ (.A1(_01074_),
    .A2(_01221_),
    .A3(_01252_),
    .B1(_01095_),
    .X(_01253_));
 sky130_fd_sc_hd__and2_1 _05979_ (.A(_01234_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__clkbuf_1 _05980_ (.A(_01254_),
    .X(\u_decod.dec0.access_size_o[0] ));
 sky130_fd_sc_hd__and2_1 _05981_ (.A(_01071_),
    .B(_01253_),
    .X(_01255_));
 sky130_fd_sc_hd__clkbuf_1 _05982_ (.A(_01255_),
    .X(\u_decod.dec0.access_size_o[1] ));
 sky130_fd_sc_hd__and4_1 _05983_ (.A(_01234_),
    .B(_01074_),
    .C(_01078_),
    .D(_01252_),
    .X(_01256_));
 sky130_fd_sc_hd__clkbuf_1 _05984_ (.A(_01256_),
    .X(\u_decod.dec0.access_size_o[2] ));
 sky130_fd_sc_hd__nand2_1 _05985_ (.A(\u_decod.rd_v_q ),
    .B(_01056_),
    .Y(_01257_));
 sky130_fd_sc_hd__inv_2 _05986_ (.A(_01257_),
    .Y(\u_decod.exe_ff_write_v_q_i ));
 sky130_fd_sc_hd__and2_1 _05987_ (.A(\u_decod.instr_unit_q[0] ),
    .B(_01056_),
    .X(_01258_));
 sky130_fd_sc_hd__buf_2 _05988_ (.A(_01258_),
    .X(_01259_));
 sky130_fd_sc_hd__buf_4 _05989_ (.A(_01259_),
    .X(_01260_));
 sky130_fd_sc_hd__nor2_1 _05990_ (.A(\u_decod.rs2_data_q[29] ),
    .B(\u_decod.rs1_data_q[29] ),
    .Y(_01261_));
 sky130_fd_sc_hd__and2_1 _05991_ (.A(\u_decod.rs2_data_q[29] ),
    .B(\u_decod.rs1_data_q[29] ),
    .X(_01262_));
 sky130_fd_sc_hd__nor2_2 _05992_ (.A(_01261_),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__and2_1 _05993_ (.A(\u_decod.rs2_data_q[28] ),
    .B(\u_decod.rs1_data_q[28] ),
    .X(_01264_));
 sky130_fd_sc_hd__nor2_1 _05994_ (.A(\u_decod.rs2_data_q[28] ),
    .B(\u_decod.rs1_data_q[28] ),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _05995_ (.A(_01264_),
    .B(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__clkbuf_4 _05996_ (.A(\u_decod.rs1_data_q[31] ),
    .X(_01267_));
 sky130_fd_sc_hd__and2_1 _05997_ (.A(\u_decod.rs2_data_q[31] ),
    .B(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_1 _05998_ (.A(\u_decod.rs2_data_q[31] ),
    .B(_01267_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _05999_ (.A(_01268_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _06000_ (.A(\u_decod.rs2_data_q[30] ),
    .B(\u_decod.rs1_data_q[30] ),
    .Y(_01271_));
 sky130_fd_sc_hd__and2_1 _06001_ (.A(\u_decod.rs2_data_q[30] ),
    .B(\u_decod.rs1_data_q[30] ),
    .X(_01272_));
 sky130_fd_sc_hd__nor2_1 _06002_ (.A(_01271_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand4_1 _06003_ (.A(_01263_),
    .B(_01266_),
    .C(_01270_),
    .D(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__or2_1 _06004_ (.A(\u_decod.rs2_data_q[25] ),
    .B(\u_decod.rs1_data_q[25] ),
    .X(_01275_));
 sky130_fd_sc_hd__nand2_1 _06005_ (.A(\u_decod.rs2_data_q[25] ),
    .B(\u_decod.rs1_data_q[25] ),
    .Y(_01276_));
 sky130_fd_sc_hd__and2_1 _06006_ (.A(_01275_),
    .B(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__nand2_2 _06007_ (.A(\u_decod.rs2_data_q[24] ),
    .B(\u_decod.rs1_data_q[24] ),
    .Y(_01278_));
 sky130_fd_sc_hd__or2_1 _06008_ (.A(\u_decod.rs2_data_q[24] ),
    .B(\u_decod.rs1_data_q[24] ),
    .X(_01279_));
 sky130_fd_sc_hd__and2_1 _06009_ (.A(_01278_),
    .B(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_1 _06010_ (.A(\u_decod.rs2_data_q[27] ),
    .B(\u_decod.rs1_data_q[27] ),
    .Y(_01281_));
 sky130_fd_sc_hd__or2_1 _06011_ (.A(\u_decod.rs2_data_q[27] ),
    .B(\u_decod.rs1_data_q[27] ),
    .X(_01282_));
 sky130_fd_sc_hd__and2_1 _06012_ (.A(_01281_),
    .B(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__or2_1 _06013_ (.A(\u_decod.rs2_data_q[26] ),
    .B(\u_decod.rs1_data_q[26] ),
    .X(_01284_));
 sky130_fd_sc_hd__nand2_1 _06014_ (.A(\u_decod.rs2_data_q[26] ),
    .B(\u_decod.rs1_data_q[26] ),
    .Y(_01285_));
 sky130_fd_sc_hd__and2_1 _06015_ (.A(_01284_),
    .B(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__nand4_1 _06016_ (.A(_01277_),
    .B(_01280_),
    .C(_01283_),
    .D(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _06017_ (.A(_01274_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__clkbuf_4 _06018_ (.A(\u_decod.rs1_data_q[15] ),
    .X(_01289_));
 sky130_fd_sc_hd__and2_2 _06019_ (.A(\u_decod.rs2_data_q[15] ),
    .B(_01289_),
    .X(_01290_));
 sky130_fd_sc_hd__nor2_1 _06020_ (.A(\u_decod.rs2_data_q[15] ),
    .B(_01289_),
    .Y(_01291_));
 sky130_fd_sc_hd__clkbuf_4 _06021_ (.A(\u_decod.rs1_data_q[14] ),
    .X(_01292_));
 sky130_fd_sc_hd__nand2_1 _06022_ (.A(\u_decod.rs2_data_q[14] ),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _06023_ (.A(_01291_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__and2_2 _06024_ (.A(\u_decod.rs2_data_q[13] ),
    .B(\u_decod.rs1_data_q[13] ),
    .X(_01295_));
 sky130_fd_sc_hd__nor2_1 _06025_ (.A(\u_decod.rs2_data_q[13] ),
    .B(\u_decod.rs1_data_q[13] ),
    .Y(_01296_));
 sky130_fd_sc_hd__clkbuf_4 _06026_ (.A(\u_decod.rs1_data_q[12] ),
    .X(_01297_));
 sky130_fd_sc_hd__nand2_1 _06027_ (.A(\u_decod.rs2_data_q[12] ),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _06028_ (.A(_01296_),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__and2_1 _06029_ (.A(\u_decod.rs2_data_q[11] ),
    .B(\u_decod.rs1_data_q[11] ),
    .X(_01300_));
 sky130_fd_sc_hd__nor2_1 _06030_ (.A(\u_decod.rs2_data_q[11] ),
    .B(\u_decod.rs1_data_q[11] ),
    .Y(_01301_));
 sky130_fd_sc_hd__clkbuf_4 _06031_ (.A(\u_decod.rs1_data_q[10] ),
    .X(_01302_));
 sky130_fd_sc_hd__nand2_1 _06032_ (.A(\u_decod.rs2_data_q[10] ),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _06033_ (.A(_01301_),
    .B(_01303_),
    .Y(_01304_));
 sky130_fd_sc_hd__and2_2 _06034_ (.A(\u_decod.rs2_data_q[9] ),
    .B(\u_decod.rs1_data_q[9] ),
    .X(_01305_));
 sky130_fd_sc_hd__nor2_1 _06035_ (.A(\u_decod.rs2_data_q[9] ),
    .B(\u_decod.rs1_data_q[9] ),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_2 _06036_ (.A(\u_decod.rs2_data_q[8] ),
    .B(\u_decod.rs1_data_q[8] ),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_1 _06037_ (.A(_01306_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _06038_ (.A(\u_decod.rs2_data_q[5] ),
    .B(\u_decod.rs1_data_q[5] ),
    .Y(_01309_));
 sky130_fd_sc_hd__nand2_1 _06039_ (.A(\u_decod.rs2_data_q[5] ),
    .B(\u_decod.rs1_data_q[5] ),
    .Y(_01310_));
 sky130_fd_sc_hd__or2b_2 _06040_ (.A(_01309_),
    .B_N(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__nor2_1 _06041_ (.A(\u_decod.rs1_data_q[3] ),
    .B(\u_decod.rs2_data_q[3] ),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _06042_ (.A(\u_decod.rs1_data_q[2] ),
    .B(\u_decod.rs2_data_q[2] ),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _06043_ (.A(\u_decod.rs1_data_q[0] ),
    .B(\u_decod.rs2_data_q[0] ),
    .Y(_01314_));
 sky130_fd_sc_hd__clkbuf_4 _06044_ (.A(\u_decod.rs2_data_q[1] ),
    .X(_01315_));
 sky130_fd_sc_hd__xnor2_2 _06045_ (.A(\u_decod.rs1_data_q[1] ),
    .B(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _06046_ (.A(\u_decod.rs1_data_q[2] ),
    .B(\u_decod.rs2_data_q[2] ),
    .Y(_01317_));
 sky130_fd_sc_hd__nand2_1 _06047_ (.A(\u_decod.rs1_data_q[1] ),
    .B(_01315_),
    .Y(_01318_));
 sky130_fd_sc_hd__o211a_1 _06048_ (.A1(_01314_),
    .A2(_01316_),
    .B1(_01317_),
    .C1(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__nand2_1 _06049_ (.A(\u_decod.rs1_data_q[3] ),
    .B(\u_decod.rs2_data_q[3] ),
    .Y(_01320_));
 sky130_fd_sc_hd__o31ai_2 _06050_ (.A1(_01312_),
    .A2(_01313_),
    .A3(_01319_),
    .B1(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__or2_1 _06051_ (.A(\u_decod.rs1_data_q[4] ),
    .B(\u_decod.rs2_data_q[4] ),
    .X(_01322_));
 sky130_fd_sc_hd__nand2_1 _06052_ (.A(\u_decod.rs1_data_q[4] ),
    .B(\u_decod.rs2_data_q[4] ),
    .Y(_01323_));
 sky130_fd_sc_hd__and2_1 _06053_ (.A(_01322_),
    .B(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__nor2_1 _06054_ (.A(\u_decod.rs2_data_q[7] ),
    .B(\u_decod.rs1_data_q[7] ),
    .Y(_01325_));
 sky130_fd_sc_hd__and2_1 _06055_ (.A(\u_decod.rs2_data_q[7] ),
    .B(\u_decod.rs1_data_q[7] ),
    .X(_01326_));
 sky130_fd_sc_hd__nor2_1 _06056_ (.A(_01325_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _06057_ (.A(\u_decod.rs2_data_q[6] ),
    .B(\u_decod.rs1_data_q[6] ),
    .Y(_01328_));
 sky130_fd_sc_hd__and2_1 _06058_ (.A(\u_decod.rs2_data_q[6] ),
    .B(\u_decod.rs1_data_q[6] ),
    .X(_01329_));
 sky130_fd_sc_hd__nor2_1 _06059_ (.A(_01328_),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__and3_1 _06060_ (.A(_01324_),
    .B(_01327_),
    .C(_01330_),
    .X(_01331_));
 sky130_fd_sc_hd__and3b_1 _06061_ (.A_N(_01311_),
    .B(_01321_),
    .C(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__a21o_1 _06062_ (.A1(_01310_),
    .A2(_01323_),
    .B1(_01309_),
    .X(_01333_));
 sky130_fd_sc_hd__nor2_1 _06063_ (.A(_01328_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__or2_1 _06064_ (.A(\u_decod.rs2_data_q[7] ),
    .B(\u_decod.rs1_data_q[7] ),
    .X(_01335_));
 sky130_fd_sc_hd__o31a_1 _06065_ (.A1(_01326_),
    .A2(_01329_),
    .A3(_01334_),
    .B1(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__nor2_1 _06066_ (.A(_01306_),
    .B(_01305_),
    .Y(_01337_));
 sky130_fd_sc_hd__inv_2 _06067_ (.A(_01307_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _06068_ (.A(\u_decod.rs2_data_q[8] ),
    .B(\u_decod.rs1_data_q[8] ),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _06069_ (.A(_01338_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__o211a_1 _06070_ (.A1(_01332_),
    .A2(_01336_),
    .B1(_01337_),
    .C1(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__nor2_1 _06071_ (.A(_01301_),
    .B(_01300_),
    .Y(_01342_));
 sky130_fd_sc_hd__and2_1 _06072_ (.A(\u_decod.rs2_data_q[10] ),
    .B(\u_decod.rs1_data_q[10] ),
    .X(_01343_));
 sky130_fd_sc_hd__nor2_1 _06073_ (.A(\u_decod.rs2_data_q[10] ),
    .B(_01302_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _06074_ (.A(_01343_),
    .B(_01344_),
    .Y(_01345_));
 sky130_fd_sc_hd__o311a_1 _06075_ (.A1(_01305_),
    .A2(_01308_),
    .A3(_01341_),
    .B1(_01342_),
    .C1(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__nor2_1 _06076_ (.A(_01296_),
    .B(_01295_),
    .Y(_01347_));
 sky130_fd_sc_hd__and2_1 _06077_ (.A(\u_decod.rs2_data_q[12] ),
    .B(_01297_),
    .X(_01348_));
 sky130_fd_sc_hd__nor2_1 _06078_ (.A(\u_decod.rs2_data_q[12] ),
    .B(_01297_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _06079_ (.A(_01348_),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__o311a_1 _06080_ (.A1(_01300_),
    .A2(_01304_),
    .A3(_01346_),
    .B1(_01347_),
    .C1(_01350_),
    .X(_01351_));
 sky130_fd_sc_hd__nor2_1 _06081_ (.A(_01291_),
    .B(_01290_),
    .Y(_01352_));
 sky130_fd_sc_hd__and2_1 _06082_ (.A(\u_decod.rs2_data_q[14] ),
    .B(_01292_),
    .X(_01353_));
 sky130_fd_sc_hd__nor2_1 _06083_ (.A(\u_decod.rs2_data_q[14] ),
    .B(_01292_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _06084_ (.A(_01353_),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__o311a_1 _06085_ (.A1(_01295_),
    .A2(_01299_),
    .A3(_01351_),
    .B1(_01352_),
    .C1(_01355_),
    .X(_01356_));
 sky130_fd_sc_hd__or3_2 _06086_ (.A(_01290_),
    .B(_01294_),
    .C(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__buf_4 _06087_ (.A(\u_decod.rs1_data_q[21] ),
    .X(_01358_));
 sky130_fd_sc_hd__nand2_1 _06088_ (.A(\u_decod.rs2_data_q[21] ),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__or2_1 _06089_ (.A(\u_decod.rs2_data_q[21] ),
    .B(_01358_),
    .X(_01360_));
 sky130_fd_sc_hd__and2_1 _06090_ (.A(_01359_),
    .B(_01360_),
    .X(_01361_));
 sky130_fd_sc_hd__inv_2 _06091_ (.A(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__clkbuf_4 _06092_ (.A(\u_decod.rs1_data_q[20] ),
    .X(_01363_));
 sky130_fd_sc_hd__and2_1 _06093_ (.A(\u_decod.rs2_data_q[20] ),
    .B(_01363_),
    .X(_01364_));
 sky130_fd_sc_hd__nor2_1 _06094_ (.A(\u_decod.rs2_data_q[20] ),
    .B(_01363_),
    .Y(_01365_));
 sky130_fd_sc_hd__or2_1 _06095_ (.A(_01364_),
    .B(_01365_),
    .X(_01366_));
 sky130_fd_sc_hd__clkbuf_4 _06096_ (.A(\u_decod.rs1_data_q[23] ),
    .X(_01367_));
 sky130_fd_sc_hd__nor2_1 _06097_ (.A(\u_decod.rs2_data_q[23] ),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__and2_1 _06098_ (.A(\u_decod.rs2_data_q[23] ),
    .B(_01367_),
    .X(_01369_));
 sky130_fd_sc_hd__or2_1 _06099_ (.A(_01368_),
    .B(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__clkbuf_4 _06100_ (.A(\u_decod.rs1_data_q[22] ),
    .X(_01371_));
 sky130_fd_sc_hd__or2_1 _06101_ (.A(\u_decod.rs2_data_q[22] ),
    .B(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__nand2_1 _06102_ (.A(\u_decod.rs2_data_q[22] ),
    .B(_01371_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _06103_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__or4_1 _06104_ (.A(_01362_),
    .B(_01366_),
    .C(_01370_),
    .D(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__clkbuf_4 _06105_ (.A(\u_decod.rs1_data_q[19] ),
    .X(_01376_));
 sky130_fd_sc_hd__or2_1 _06106_ (.A(\u_decod.rs2_data_q[19] ),
    .B(_01376_),
    .X(_01377_));
 sky130_fd_sc_hd__nand2_1 _06107_ (.A(\u_decod.rs2_data_q[19] ),
    .B(_01376_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _06108_ (.A(_01377_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__clkbuf_4 _06109_ (.A(\u_decod.rs1_data_q[17] ),
    .X(_01380_));
 sky130_fd_sc_hd__nand2_1 _06110_ (.A(\u_decod.rs2_data_q[17] ),
    .B(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__or2_1 _06111_ (.A(\u_decod.rs2_data_q[17] ),
    .B(_01380_),
    .X(_01382_));
 sky130_fd_sc_hd__nand2_1 _06112_ (.A(_01381_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__clkbuf_4 _06113_ (.A(\u_decod.rs1_data_q[18] ),
    .X(_01384_));
 sky130_fd_sc_hd__or2_1 _06114_ (.A(\u_decod.rs2_data_q[18] ),
    .B(_01384_),
    .X(_01385_));
 sky130_fd_sc_hd__nand2_1 _06115_ (.A(\u_decod.rs2_data_q[18] ),
    .B(_01384_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _06116_ (.A(_01385_),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__clkbuf_4 _06117_ (.A(\u_decod.rs1_data_q[16] ),
    .X(_01388_));
 sky130_fd_sc_hd__and2_1 _06118_ (.A(\u_decod.rs2_data_q[16] ),
    .B(_01388_),
    .X(_01389_));
 sky130_fd_sc_hd__nor2_1 _06119_ (.A(\u_decod.rs2_data_q[16] ),
    .B(_01388_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_2 _06120_ (.A(_01389_),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__or4b_1 _06121_ (.A(_01379_),
    .B(_01383_),
    .C(_01387_),
    .D_N(_01391_),
    .X(_01392_));
 sky130_fd_sc_hd__nor2_1 _06122_ (.A(_01375_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand3_1 _06123_ (.A(_01288_),
    .B(_01357_),
    .C(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _06124_ (.A(\u_decod.rs2_data_q[20] ),
    .B(_01363_),
    .Y(_01395_));
 sky130_fd_sc_hd__nor2_1 _06125_ (.A(\u_decod.rs2_data_q[21] ),
    .B(_01358_),
    .Y(_01396_));
 sky130_fd_sc_hd__a21oi_1 _06126_ (.A1(_01359_),
    .A2(_01395_),
    .B1(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__and2_1 _06127_ (.A(\u_decod.rs2_data_q[22] ),
    .B(_01371_),
    .X(_01398_));
 sky130_fd_sc_hd__o221a_1 _06128_ (.A1(\u_decod.rs2_data_q[23] ),
    .A2(_01367_),
    .B1(_01397_),
    .B2(_01398_),
    .C1(_01372_),
    .X(_01399_));
 sky130_fd_sc_hd__nand2_2 _06129_ (.A(\u_decod.rs2_data_q[16] ),
    .B(_01388_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _06130_ (.A(\u_decod.rs2_data_q[17] ),
    .B(_01380_),
    .Y(_01401_));
 sky130_fd_sc_hd__a21oi_1 _06131_ (.A1(_01381_),
    .A2(_01400_),
    .B1(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__and2_1 _06132_ (.A(\u_decod.rs2_data_q[18] ),
    .B(_01384_),
    .X(_01403_));
 sky130_fd_sc_hd__a221o_1 _06133_ (.A1(\u_decod.rs2_data_q[19] ),
    .A2(_01376_),
    .B1(_01385_),
    .B2(_01402_),
    .C1(_01403_),
    .X(_01404_));
 sky130_fd_sc_hd__nand2_2 _06134_ (.A(_01377_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _06135_ (.A(_01375_),
    .B(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__or3_2 _06136_ (.A(_01369_),
    .B(_01399_),
    .C(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__nand2_1 _06137_ (.A(_01288_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__and2_1 _06138_ (.A(\u_decod.rs2_data_q[26] ),
    .B(\u_decod.rs1_data_q[26] ),
    .X(_01409_));
 sky130_fd_sc_hd__nor2_1 _06139_ (.A(\u_decod.rs2_data_q[25] ),
    .B(\u_decod.rs1_data_q[25] ),
    .Y(_01410_));
 sky130_fd_sc_hd__a21oi_1 _06140_ (.A1(_01276_),
    .A2(_01278_),
    .B1(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__o21a_1 _06141_ (.A1(_01409_),
    .A2(_01411_),
    .B1(_01282_),
    .X(_01412_));
 sky130_fd_sc_hd__a21boi_1 _06142_ (.A1(_01284_),
    .A2(_01412_),
    .B1_N(_01281_),
    .Y(_01413_));
 sky130_fd_sc_hd__or2_1 _06143_ (.A(\u_decod.rs2_data_q[29] ),
    .B(\u_decod.rs1_data_q[29] ),
    .X(_01414_));
 sky130_fd_sc_hd__o21a_1 _06144_ (.A1(_01262_),
    .A2(_01264_),
    .B1(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__o21bai_1 _06145_ (.A1(_01272_),
    .A2(_01415_),
    .B1_N(_01269_),
    .Y(_01416_));
 sky130_fd_sc_hd__o21ba_1 _06146_ (.A1(_01271_),
    .A2(_01416_),
    .B1_N(_01268_),
    .X(_01417_));
 sky130_fd_sc_hd__o21a_1 _06147_ (.A1(_01274_),
    .A2(_01413_),
    .B1(_01417_),
    .X(_01418_));
 sky130_fd_sc_hd__xnor2_4 _06148_ (.A(\u_decod.rs2_data_q[32] ),
    .B(\u_decod.rs1_data_q[32] ),
    .Y(_01419_));
 sky130_fd_sc_hd__a31o_1 _06149_ (.A1(_01394_),
    .A2(_01408_),
    .A3(_01418_),
    .B1(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__nand4_2 _06150_ (.A(_01394_),
    .B(_01408_),
    .C(_01418_),
    .D(_01419_),
    .Y(_01421_));
 sky130_fd_sc_hd__buf_2 _06151_ (.A(\u_decod.rs2_data_q[0] ),
    .X(_01422_));
 sky130_fd_sc_hd__buf_2 _06152_ (.A(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__buf_2 _06153_ (.A(_01423_),
    .X(_01424_));
 sky130_fd_sc_hd__buf_2 _06154_ (.A(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__or2_1 _06155_ (.A(_01061_),
    .B(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__clkbuf_4 _06156_ (.A(_01056_),
    .X(_01427_));
 sky130_fd_sc_hd__and3_1 _06157_ (.A(\u_decod.instr_unit_q[0] ),
    .B(\u_decod.instr_operation_q[1] ),
    .C(_01427_),
    .X(_01428_));
 sky130_fd_sc_hd__clkbuf_4 _06158_ (.A(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__buf_4 _06159_ (.A(\u_decod.instr_operation_q[2] ),
    .X(_01430_));
 sky130_fd_sc_hd__and3_2 _06160_ (.A(\u_decod.instr_unit_q[0] ),
    .B(_01430_),
    .C(_01427_),
    .X(_01431_));
 sky130_fd_sc_hd__clkbuf_4 _06161_ (.A(_01431_),
    .X(_01432_));
 sky130_fd_sc_hd__and3_1 _06162_ (.A(\u_decod.instr_unit_q[0] ),
    .B(\u_decod.instr_operation_q[3] ),
    .C(_01056_),
    .X(_01433_));
 sky130_fd_sc_hd__clkbuf_2 _06163_ (.A(_01433_),
    .X(_01434_));
 sky130_fd_sc_hd__clkbuf_4 _06164_ (.A(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__and3_2 _06165_ (.A(\u_decod.instr_unit_q[0] ),
    .B(\u_decod.instr_operation_q[0] ),
    .C(_01427_),
    .X(_01436_));
 sky130_fd_sc_hd__clkbuf_4 _06166_ (.A(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__o21a_1 _06167_ (.A1(_01435_),
    .A2(_01437_),
    .B1(_01314_),
    .X(_01438_));
 sky130_fd_sc_hd__a311o_1 _06168_ (.A1(_01061_),
    .A2(_01425_),
    .A3(_01429_),
    .B1(_01432_),
    .C1(_01438_),
    .X(_01439_));
 sky130_fd_sc_hd__a32o_1 _06169_ (.A1(\u_decod.instr_operation_q[4] ),
    .A2(_01420_),
    .A3(_01421_),
    .B1(_01426_),
    .B2(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__o211a_4 _06170_ (.A1(\u_decod.instr_operation_q[1] ),
    .A2(_01430_),
    .B1(\u_decod.instr_unit_q[1] ),
    .C1(_01427_),
    .X(_01441_));
 sky130_fd_sc_hd__buf_2 _06171_ (.A(_01441_),
    .X(_01442_));
 sky130_fd_sc_hd__buf_2 _06172_ (.A(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__clkbuf_4 _06173_ (.A(\u_decod.rs2_data_q[3] ),
    .X(_01444_));
 sky130_fd_sc_hd__buf_2 _06174_ (.A(\u_decod.rs2_data_q[4] ),
    .X(_01445_));
 sky130_fd_sc_hd__clkbuf_4 _06175_ (.A(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__buf_2 _06176_ (.A(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__mux4_1 _06177_ (.A0(\u_decod.rs1_data_q[3] ),
    .A1(\u_decod.rs1_data_q[11] ),
    .A2(_01376_),
    .A3(\u_decod.rs1_data_q[27] ),
    .S0(_01444_),
    .S1(_01447_),
    .X(_01448_));
 sky130_fd_sc_hd__mux4_1 _06178_ (.A0(\u_decod.rs1_data_q[7] ),
    .A1(_01289_),
    .A2(_01367_),
    .A3(_01267_),
    .S0(_01444_),
    .S1(_01447_),
    .X(_01449_));
 sky130_fd_sc_hd__clkbuf_4 _06179_ (.A(\u_decod.rs2_data_q[2] ),
    .X(_01450_));
 sky130_fd_sc_hd__clkbuf_4 _06180_ (.A(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _06181_ (.A0(_01448_),
    .A1(_01449_),
    .S(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__mux4_1 _06182_ (.A0(\u_decod.rs1_data_q[5] ),
    .A1(\u_decod.rs1_data_q[13] ),
    .A2(_01358_),
    .A3(\u_decod.rs1_data_q[29] ),
    .S0(_01444_),
    .S1(_01447_),
    .X(_01453_));
 sky130_fd_sc_hd__buf_2 _06183_ (.A(_01445_),
    .X(_01454_));
 sky130_fd_sc_hd__clkbuf_4 _06184_ (.A(\u_decod.rs2_data_q[3] ),
    .X(_01455_));
 sky130_fd_sc_hd__mux4_1 _06185_ (.A0(\u_decod.rs1_data_q[1] ),
    .A1(_01380_),
    .A2(\u_decod.rs1_data_q[9] ),
    .A3(\u_decod.rs1_data_q[25] ),
    .S0(_01454_),
    .S1(_01455_),
    .X(_01456_));
 sky130_fd_sc_hd__inv_2 _06186_ (.A(_01450_),
    .Y(_01457_));
 sky130_fd_sc_hd__clkbuf_4 _06187_ (.A(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _06188_ (.A0(_01453_),
    .A1(_01456_),
    .S(_01458_),
    .X(_01459_));
 sky130_fd_sc_hd__clkbuf_4 _06189_ (.A(_01444_),
    .X(_01460_));
 sky130_fd_sc_hd__buf_2 _06190_ (.A(_01447_),
    .X(_01461_));
 sky130_fd_sc_hd__mux4_1 _06191_ (.A0(\u_decod.rs1_data_q[2] ),
    .A1(_01302_),
    .A2(_01384_),
    .A3(\u_decod.rs1_data_q[26] ),
    .S0(_01460_),
    .S1(_01461_),
    .X(_01462_));
 sky130_fd_sc_hd__mux4_1 _06192_ (.A0(\u_decod.rs1_data_q[6] ),
    .A1(_01292_),
    .A2(_01371_),
    .A3(\u_decod.rs1_data_q[30] ),
    .S0(_01444_),
    .S1(_01447_),
    .X(_01463_));
 sky130_fd_sc_hd__clkbuf_4 _06193_ (.A(_01451_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _06194_ (.A0(_01462_),
    .A1(_01463_),
    .S(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__clkbuf_4 _06195_ (.A(_01461_),
    .X(_01466_));
 sky130_fd_sc_hd__clkbuf_4 _06196_ (.A(_01455_),
    .X(_01467_));
 sky130_fd_sc_hd__clkbuf_4 _06197_ (.A(_01467_),
    .X(_01468_));
 sky130_fd_sc_hd__clkbuf_4 _06198_ (.A(_01468_),
    .X(_01469_));
 sky130_fd_sc_hd__mux4_1 _06199_ (.A0(_01061_),
    .A1(_01388_),
    .A2(\u_decod.rs1_data_q[8] ),
    .A3(\u_decod.rs1_data_q[24] ),
    .S0(_01466_),
    .S1(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__mux4_1 _06200_ (.A0(\u_decod.rs1_data_q[4] ),
    .A1(_01297_),
    .A2(_01363_),
    .A3(\u_decod.rs1_data_q[28] ),
    .S0(_01460_),
    .S1(_01461_),
    .X(_01471_));
 sky130_fd_sc_hd__buf_2 _06201_ (.A(_01451_),
    .X(_01472_));
 sky130_fd_sc_hd__mux2_1 _06202_ (.A0(_01470_),
    .A1(_01471_),
    .S(_01472_),
    .X(_01473_));
 sky130_fd_sc_hd__inv_2 _06203_ (.A(_01315_),
    .Y(_01474_));
 sky130_fd_sc_hd__clkbuf_4 _06204_ (.A(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__clkbuf_4 _06205_ (.A(_01475_),
    .X(_01476_));
 sky130_fd_sc_hd__clkbuf_4 _06206_ (.A(_01476_),
    .X(_01477_));
 sky130_fd_sc_hd__inv_2 _06207_ (.A(\u_decod.rs2_data_q[0] ),
    .Y(_01478_));
 sky130_fd_sc_hd__buf_2 _06208_ (.A(_01478_),
    .X(_01479_));
 sky130_fd_sc_hd__clkbuf_4 _06209_ (.A(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__clkbuf_4 _06210_ (.A(_01480_),
    .X(_01481_));
 sky130_fd_sc_hd__mux4_1 _06211_ (.A0(_01452_),
    .A1(_01459_),
    .A2(_01465_),
    .A3(_01473_),
    .S0(_01477_),
    .S1(_01481_),
    .X(_01482_));
 sky130_fd_sc_hd__and2_1 _06212_ (.A(\u_decod.instr_unit_q[2] ),
    .B(_01056_),
    .X(_01483_));
 sky130_fd_sc_hd__clkbuf_2 _06213_ (.A(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__buf_4 _06214_ (.A(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__or2_1 _06215_ (.A(net98),
    .B(net99),
    .X(_01486_));
 sky130_fd_sc_hd__a31o_2 _06216_ (.A1(_01064_),
    .A2(_01067_),
    .A3(_01486_),
    .B1(net100),
    .X(_01487_));
 sky130_fd_sc_hd__and3_2 _06217_ (.A(net112),
    .B(_01066_),
    .C(_01486_),
    .X(_01488_));
 sky130_fd_sc_hd__and3b_2 _06218_ (.A_N(_01063_),
    .B(net101),
    .C(net98),
    .X(_01489_));
 sky130_fd_sc_hd__and3_2 _06219_ (.A(net98),
    .B(_01063_),
    .C(net101),
    .X(_01490_));
 sky130_fd_sc_hd__a22o_1 _06220_ (.A1(net63),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net49),
    .X(_01491_));
 sky130_fd_sc_hd__a221o_1 _06221_ (.A1(net33),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net40),
    .C1(_01491_),
    .X(_01492_));
 sky130_fd_sc_hd__buf_2 _06222_ (.A(_01315_),
    .X(_01493_));
 sky130_fd_sc_hd__a21bo_1 _06223_ (.A1(\u_decod.rs1_data_q[31] ),
    .A2(\u_decod.instr_operation_q[2] ),
    .B1_N(_01445_),
    .X(_01494_));
 sky130_fd_sc_hd__o21a_1 _06224_ (.A1(_01061_),
    .A2(_01445_),
    .B1(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__nand2_2 _06225_ (.A(_01267_),
    .B(_01430_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_2 _06226_ (.A(\u_decod.rs2_data_q[3] ),
    .B(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__buf_2 _06227_ (.A(_01497_),
    .X(_01498_));
 sky130_fd_sc_hd__o21a_1 _06228_ (.A1(_01460_),
    .A2(_01495_),
    .B1(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__nand2_2 _06229_ (.A(_01450_),
    .B(_01496_),
    .Y(_01500_));
 sky130_fd_sc_hd__o21a_1 _06230_ (.A1(_01451_),
    .A2(_01499_),
    .B1(_01500_),
    .X(_01501_));
 sky130_fd_sc_hd__nand2_1 _06231_ (.A(_01315_),
    .B(_01496_),
    .Y(_01502_));
 sky130_fd_sc_hd__o21a_1 _06232_ (.A1(_01493_),
    .A2(_01501_),
    .B1(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__and3_1 _06233_ (.A(\u_decod.instr_operation_q[0] ),
    .B(\u_decod.instr_unit_q[1] ),
    .C(_01427_),
    .X(_01504_));
 sky130_fd_sc_hd__buf_2 _06234_ (.A(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__clkbuf_4 _06235_ (.A(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__nand2_1 _06236_ (.A(_01424_),
    .B(_01496_),
    .Y(_01507_));
 sky130_fd_sc_hd__o211a_1 _06237_ (.A1(_01424_),
    .A2(_01503_),
    .B1(_01506_),
    .C1(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__a221o_1 _06238_ (.A1(\u_decod.pc_q_o[0] ),
    .A2(_01485_),
    .B1(_01492_),
    .B2(_01059_),
    .C1(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__a21o_1 _06239_ (.A1(_01443_),
    .A2(_01482_),
    .B1(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__a21oi_2 _06240_ (.A1(_01260_),
    .A2(_01440_),
    .B1(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__inv_2 _06241_ (.A(_01511_),
    .Y(\u_decod.exe_ff_res_data_i[0] ));
 sky130_fd_sc_hd__inv_2 _06242_ (.A(\u_decod.dec0.instr_i[24] ),
    .Y(_01512_));
 sky130_fd_sc_hd__clkbuf_2 _06243_ (.A(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__nor2_1 _06244_ (.A(\u_decod.dec0.instr_i[20] ),
    .B(\u_decod.dec0.instr_i[21] ),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_2 _06245_ (.A(\u_decod.dec0.instr_i[22] ),
    .B(\u_decod.dec0.instr_i[23] ),
    .Y(_01515_));
 sky130_fd_sc_hd__and3_4 _06246_ (.A(_01513_),
    .B(_01514_),
    .C(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__a211oi_4 _06247_ (.A1(\u_decod.dec0.instr_i[6] ),
    .A2(\u_decod.dec0.instr_i[4] ),
    .B1(_01225_),
    .C1(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__inv_2 _06248_ (.A(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__xor2_1 _06249_ (.A(\u_decod.dec0.instr_i[23] ),
    .B(\u_decod.exe_ff_rd_adr_q_i[3] ),
    .X(_01519_));
 sky130_fd_sc_hd__inv_2 _06250_ (.A(\u_decod.dec0.instr_i[20] ),
    .Y(_01520_));
 sky130_fd_sc_hd__inv_2 _06251_ (.A(\u_decod.exe_ff_rd_adr_q_i[1] ),
    .Y(_01521_));
 sky130_fd_sc_hd__inv_2 _06252_ (.A(\u_decod.dec0.instr_i[22] ),
    .Y(_01522_));
 sky130_fd_sc_hd__a22o_1 _06253_ (.A1(\u_decod.dec0.instr_i[21] ),
    .A2(_01521_),
    .B1(\u_decod.exe_ff_rd_adr_q_i[2] ),
    .B2(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__a221o_1 _06254_ (.A1(_01520_),
    .A2(\u_decod.exe_ff_rd_adr_q_i[0] ),
    .B1(\u_decod.exe_ff_rd_adr_q_i[4] ),
    .B2(_01512_),
    .C1(_01523_),
    .X(_01524_));
 sky130_fd_sc_hd__o22a_1 _06255_ (.A1(_01520_),
    .A2(\u_decod.exe_ff_rd_adr_q_i[0] ),
    .B1(\u_decod.exe_ff_rd_adr_q_i[2] ),
    .B2(_01522_),
    .X(_01525_));
 sky130_fd_sc_hd__o221ai_1 _06256_ (.A1(\u_decod.dec0.instr_i[21] ),
    .A2(_01521_),
    .B1(\u_decod.exe_ff_rd_adr_q_i[4] ),
    .B2(_01513_),
    .C1(_01525_),
    .Y(_01526_));
 sky130_fd_sc_hd__or4_2 _06257_ (.A(_01257_),
    .B(_01519_),
    .C(_01524_),
    .D(_01526_),
    .X(_01527_));
 sky130_fd_sc_hd__or2_4 _06258_ (.A(_01518_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__a21o_1 _06259_ (.A1(_01087_),
    .A2(_01199_),
    .B1(\u_decod.dec0.jalr ),
    .X(_01529_));
 sky130_fd_sc_hd__clkbuf_4 _06260_ (.A(_01529_),
    .X(_01530_));
 sky130_fd_sc_hd__buf_2 _06261_ (.A(\u_decod.rf_ff_rd_adr_q_i[2] ),
    .X(_01531_));
 sky130_fd_sc_hd__inv_2 _06262_ (.A(\u_decod.rf_ff_rd_adr_q_i[2] ),
    .Y(_01532_));
 sky130_fd_sc_hd__o22a_1 _06263_ (.A1(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .A2(_01520_),
    .B1(\u_decod.dec0.instr_i[22] ),
    .B2(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__inv_2 _06264_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .Y(_01534_));
 sky130_fd_sc_hd__inv_2 _06265_ (.A(\u_decod.rf_ff_rd_adr_q_i[3] ),
    .Y(_01535_));
 sky130_fd_sc_hd__buf_2 _06266_ (.A(\u_decod.rf_ff_rd_adr_q_i[3] ),
    .X(_01536_));
 sky130_fd_sc_hd__inv_2 _06267_ (.A(\u_decod.dec0.instr_i[23] ),
    .Y(_01537_));
 sky130_fd_sc_hd__buf_2 _06268_ (.A(\u_decod.dec0.instr_i[24] ),
    .X(_01538_));
 sky130_fd_sc_hd__inv_2 _06269_ (.A(\u_decod.rf_ff_rd_adr_q_i[4] ),
    .Y(_01539_));
 sky130_fd_sc_hd__o22a_1 _06270_ (.A1(_01536_),
    .A2(_01537_),
    .B1(_01538_),
    .B2(_01539_),
    .X(_01540_));
 sky130_fd_sc_hd__o221a_1 _06271_ (.A1(_01534_),
    .A2(\u_decod.dec0.instr_i[20] ),
    .B1(\u_decod.dec0.instr_i[23] ),
    .B2(_01535_),
    .C1(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__inv_2 _06272_ (.A(\u_decod.rf_ff_rd_adr_q_i[1] ),
    .Y(_01542_));
 sky130_fd_sc_hd__o22a_1 _06273_ (.A1(_01542_),
    .A2(\u_decod.dec0.instr_i[21] ),
    .B1(_01512_),
    .B2(\u_decod.rf_ff_rd_adr_q_i[4] ),
    .X(_01543_));
 sky130_fd_sc_hd__or2b_1 _06274_ (.A(\u_decod.flush_v ),
    .B_N(\u_decod.rf_write_v_q_i ),
    .X(_01544_));
 sky130_fd_sc_hd__a21oi_1 _06275_ (.A1(_01542_),
    .A2(\u_decod.dec0.instr_i[21] ),
    .B1(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__and3_1 _06276_ (.A(_01541_),
    .B(_01543_),
    .C(_01545_),
    .X(_01546_));
 sky130_fd_sc_hd__o211a_1 _06277_ (.A1(_01531_),
    .A2(_01522_),
    .B1(_01533_),
    .C1(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__and3_2 _06278_ (.A(_01517_),
    .B(_01527_),
    .C(_01547_),
    .X(_01548_));
 sky130_fd_sc_hd__buf_2 _06279_ (.A(_01548_),
    .X(_01549_));
 sky130_fd_sc_hd__clkbuf_4 _06280_ (.A(_01549_),
    .X(_01550_));
 sky130_fd_sc_hd__nor2_1 _06281_ (.A(_01522_),
    .B(\u_decod.dec0.instr_i[23] ),
    .Y(_01551_));
 sky130_fd_sc_hd__inv_2 _06282_ (.A(\u_decod.dec0.instr_i[21] ),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _06283_ (.A(\u_decod.dec0.instr_i[20] ),
    .B(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__and3_2 _06284_ (.A(_01512_),
    .B(_01551_),
    .C(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__clkbuf_8 _06285_ (.A(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__buf_4 _06286_ (.A(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__clkbuf_8 _06287_ (.A(_01556_),
    .X(_01557_));
 sky130_fd_sc_hd__nor2_1 _06288_ (.A(_01520_),
    .B(_01552_),
    .Y(_01558_));
 sky130_fd_sc_hd__and3_2 _06289_ (.A(_01512_),
    .B(_01551_),
    .C(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__clkbuf_8 _06290_ (.A(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__clkbuf_8 _06291_ (.A(_01560_),
    .X(_01561_));
 sky130_fd_sc_hd__clkbuf_8 _06292_ (.A(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__and3_2 _06293_ (.A(_01538_),
    .B(_01514_),
    .C(_01515_),
    .X(_01563_));
 sky130_fd_sc_hd__clkbuf_8 _06294_ (.A(_01563_),
    .X(_01564_));
 sky130_fd_sc_hd__clkbuf_8 _06295_ (.A(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _06296_ (.A(_01520_),
    .B(\u_decod.dec0.instr_i[21] ),
    .Y(_01566_));
 sky130_fd_sc_hd__and3_2 _06297_ (.A(_01513_),
    .B(_01566_),
    .C(_01551_),
    .X(_01567_));
 sky130_fd_sc_hd__clkbuf_8 _06298_ (.A(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__buf_4 _06299_ (.A(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__a22o_1 _06300_ (.A1(\u_rf.reg16_q[0] ),
    .A2(_01565_),
    .B1(_01569_),
    .B2(\u_rf.reg5_q[0] ),
    .X(_01570_));
 sky130_fd_sc_hd__a221o_1 _06301_ (.A1(\u_rf.reg6_q[0] ),
    .A2(_01557_),
    .B1(_01562_),
    .B2(\u_rf.reg7_q[0] ),
    .C1(_01570_),
    .X(_01571_));
 sky130_fd_sc_hd__buf_2 _06302_ (.A(_01538_),
    .X(_01572_));
 sky130_fd_sc_hd__nor2_1 _06303_ (.A(\u_decod.dec0.instr_i[22] ),
    .B(_01537_),
    .Y(_01573_));
 sky130_fd_sc_hd__and3_2 _06304_ (.A(_01572_),
    .B(_01566_),
    .C(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__clkbuf_8 _06305_ (.A(_01574_),
    .X(_01575_));
 sky130_fd_sc_hd__buf_6 _06306_ (.A(_01575_),
    .X(_01576_));
 sky130_fd_sc_hd__nor2_1 _06307_ (.A(_01522_),
    .B(_01537_),
    .Y(_01577_));
 sky130_fd_sc_hd__and3_2 _06308_ (.A(_01538_),
    .B(_01553_),
    .C(_01577_),
    .X(_01578_));
 sky130_fd_sc_hd__buf_6 _06309_ (.A(_01578_),
    .X(_01579_));
 sky130_fd_sc_hd__buf_6 _06310_ (.A(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__buf_6 _06311_ (.A(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__and3_2 _06312_ (.A(_01512_),
    .B(_01558_),
    .C(_01573_),
    .X(_01582_));
 sky130_fd_sc_hd__clkbuf_8 _06313_ (.A(_01582_),
    .X(_01583_));
 sky130_fd_sc_hd__buf_4 _06314_ (.A(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__and3_2 _06315_ (.A(_01513_),
    .B(_01515_),
    .C(_01566_),
    .X(_01585_));
 sky130_fd_sc_hd__clkbuf_8 _06316_ (.A(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__buf_4 _06317_ (.A(_01586_),
    .X(_01587_));
 sky130_fd_sc_hd__a22o_1 _06318_ (.A1(\u_rf.reg11_q[0] ),
    .A2(_01584_),
    .B1(_01587_),
    .B2(\u_rf.reg1_q[0] ),
    .X(_01588_));
 sky130_fd_sc_hd__a221o_1 _06319_ (.A1(\u_rf.reg25_q[0] ),
    .A2(_01576_),
    .B1(_01581_),
    .B2(\u_rf.reg30_q[0] ),
    .C1(_01588_),
    .X(_01589_));
 sky130_fd_sc_hd__and3_2 _06320_ (.A(_01572_),
    .B(_01515_),
    .C(_01553_),
    .X(_01590_));
 sky130_fd_sc_hd__clkbuf_8 _06321_ (.A(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__clkbuf_8 _06322_ (.A(_01591_),
    .X(_01592_));
 sky130_fd_sc_hd__and3_2 _06323_ (.A(_01572_),
    .B(_01515_),
    .C(_01558_),
    .X(_01593_));
 sky130_fd_sc_hd__clkbuf_8 _06324_ (.A(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__buf_4 _06325_ (.A(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__and3_2 _06326_ (.A(_01513_),
    .B(_01566_),
    .C(_01577_),
    .X(_01596_));
 sky130_fd_sc_hd__clkbuf_8 _06327_ (.A(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__clkbuf_8 _06328_ (.A(_01597_),
    .X(_01598_));
 sky130_fd_sc_hd__and3_2 _06329_ (.A(_01513_),
    .B(_01558_),
    .C(_01577_),
    .X(_01599_));
 sky130_fd_sc_hd__clkbuf_8 _06330_ (.A(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__buf_6 _06331_ (.A(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__a22o_1 _06332_ (.A1(\u_rf.reg13_q[0] ),
    .A2(_01598_),
    .B1(_01601_),
    .B2(\u_rf.reg15_q[0] ),
    .X(_01602_));
 sky130_fd_sc_hd__a221o_1 _06333_ (.A1(\u_rf.reg18_q[0] ),
    .A2(_01592_),
    .B1(_01595_),
    .B2(\u_rf.reg19_q[0] ),
    .C1(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__and3_2 _06334_ (.A(_01512_),
    .B(_01515_),
    .C(_01558_),
    .X(_01604_));
 sky130_fd_sc_hd__clkbuf_8 _06335_ (.A(_01604_),
    .X(_01605_));
 sky130_fd_sc_hd__clkbuf_8 _06336_ (.A(_01605_),
    .X(_01606_));
 sky130_fd_sc_hd__and3_2 _06337_ (.A(_01513_),
    .B(_01514_),
    .C(_01577_),
    .X(_01607_));
 sky130_fd_sc_hd__clkbuf_8 _06338_ (.A(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__buf_4 _06339_ (.A(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__clkbuf_8 _06340_ (.A(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__and3_2 _06341_ (.A(_01572_),
    .B(_01551_),
    .C(_01558_),
    .X(_01611_));
 sky130_fd_sc_hd__buf_6 _06342_ (.A(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__clkbuf_8 _06343_ (.A(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__and3_2 _06344_ (.A(_01538_),
    .B(_01558_),
    .C(_01577_),
    .X(_01614_));
 sky130_fd_sc_hd__clkbuf_8 _06345_ (.A(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__buf_4 _06346_ (.A(_01615_),
    .X(_01616_));
 sky130_fd_sc_hd__a22o_1 _06347_ (.A1(\u_rf.reg23_q[0] ),
    .A2(_01613_),
    .B1(_01616_),
    .B2(\u_rf.reg31_q[0] ),
    .X(_01617_));
 sky130_fd_sc_hd__a221o_1 _06348_ (.A1(\u_rf.reg3_q[0] ),
    .A2(_01606_),
    .B1(_01610_),
    .B2(\u_rf.reg12_q[0] ),
    .C1(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__or4_1 _06349_ (.A(_01571_),
    .B(_01589_),
    .C(_01603_),
    .D(_01618_),
    .X(_01619_));
 sky130_fd_sc_hd__and3_2 _06350_ (.A(_01572_),
    .B(_01514_),
    .C(_01573_),
    .X(_01620_));
 sky130_fd_sc_hd__buf_6 _06351_ (.A(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__clkbuf_8 _06352_ (.A(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__and3_2 _06353_ (.A(_01538_),
    .B(_01514_),
    .C(_01577_),
    .X(_01623_));
 sky130_fd_sc_hd__clkbuf_8 _06354_ (.A(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__clkbuf_8 _06355_ (.A(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__and3_2 _06356_ (.A(_01572_),
    .B(_01566_),
    .C(_01577_),
    .X(_01626_));
 sky130_fd_sc_hd__clkbuf_8 _06357_ (.A(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__buf_4 _06358_ (.A(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__and3_2 _06359_ (.A(_01538_),
    .B(_01515_),
    .C(_01566_),
    .X(_01629_));
 sky130_fd_sc_hd__clkbuf_8 _06360_ (.A(_01629_),
    .X(_01630_));
 sky130_fd_sc_hd__clkbuf_8 _06361_ (.A(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__a22o_1 _06362_ (.A1(\u_rf.reg29_q[0] ),
    .A2(_01628_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[0] ),
    .X(_01632_));
 sky130_fd_sc_hd__a221o_1 _06363_ (.A1(\u_rf.reg24_q[0] ),
    .A2(_01622_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[0] ),
    .C1(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__and3_2 _06364_ (.A(_01513_),
    .B(_01566_),
    .C(_01573_),
    .X(_01634_));
 sky130_fd_sc_hd__clkbuf_8 _06365_ (.A(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__clkbuf_8 _06366_ (.A(_01635_),
    .X(_01636_));
 sky130_fd_sc_hd__and3_2 _06367_ (.A(_01572_),
    .B(_01566_),
    .C(_01551_),
    .X(_01637_));
 sky130_fd_sc_hd__buf_6 _06368_ (.A(_01637_),
    .X(_01638_));
 sky130_fd_sc_hd__clkbuf_8 _06369_ (.A(_01638_),
    .X(_01639_));
 sky130_fd_sc_hd__and3_2 _06370_ (.A(_01538_),
    .B(_01553_),
    .C(_01573_),
    .X(_01640_));
 sky130_fd_sc_hd__clkbuf_8 _06371_ (.A(_01640_),
    .X(_01641_));
 sky130_fd_sc_hd__clkbuf_8 _06372_ (.A(_01641_),
    .X(_01642_));
 sky130_fd_sc_hd__and3_2 _06373_ (.A(_01538_),
    .B(_01514_),
    .C(_01551_),
    .X(_01643_));
 sky130_fd_sc_hd__clkbuf_8 _06374_ (.A(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__clkbuf_8 _06375_ (.A(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__a22o_1 _06376_ (.A1(\u_rf.reg26_q[0] ),
    .A2(_01642_),
    .B1(_01645_),
    .B2(\u_rf.reg20_q[0] ),
    .X(_01646_));
 sky130_fd_sc_hd__a221o_1 _06377_ (.A1(\u_rf.reg9_q[0] ),
    .A2(_01636_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[0] ),
    .C1(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__and3_2 _06378_ (.A(_01512_),
    .B(_01514_),
    .C(_01551_),
    .X(_01648_));
 sky130_fd_sc_hd__clkbuf_8 _06379_ (.A(_01648_),
    .X(_01649_));
 sky130_fd_sc_hd__clkbuf_8 _06380_ (.A(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__and3_2 _06381_ (.A(_01572_),
    .B(_01551_),
    .C(_01553_),
    .X(_01651_));
 sky130_fd_sc_hd__clkbuf_8 _06382_ (.A(_01651_),
    .X(_01652_));
 sky130_fd_sc_hd__clkbuf_8 _06383_ (.A(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__clkbuf_8 _06384_ (.A(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__and3_2 _06385_ (.A(_01513_),
    .B(_01553_),
    .C(_01573_),
    .X(_01655_));
 sky130_fd_sc_hd__clkbuf_8 _06386_ (.A(_01655_),
    .X(_01656_));
 sky130_fd_sc_hd__and3_2 _06387_ (.A(_01512_),
    .B(_01553_),
    .C(_01577_),
    .X(_01657_));
 sky130_fd_sc_hd__clkbuf_8 _06388_ (.A(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__buf_4 _06389_ (.A(_01658_),
    .X(_01659_));
 sky130_fd_sc_hd__a22o_1 _06390_ (.A1(\u_rf.reg10_q[0] ),
    .A2(_01656_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[0] ),
    .X(_01660_));
 sky130_fd_sc_hd__a221o_1 _06391_ (.A1(\u_rf.reg4_q[0] ),
    .A2(_01650_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[0] ),
    .C1(_01660_),
    .X(_01661_));
 sky130_fd_sc_hd__clkbuf_8 _06392_ (.A(_01516_),
    .X(_01662_));
 sky130_fd_sc_hd__clkbuf_8 _06393_ (.A(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__clkbuf_8 _06394_ (.A(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__and3_2 _06395_ (.A(_01512_),
    .B(_01514_),
    .C(_01573_),
    .X(_01665_));
 sky130_fd_sc_hd__clkbuf_8 _06396_ (.A(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__clkbuf_8 _06397_ (.A(_01666_),
    .X(_01667_));
 sky130_fd_sc_hd__clkbuf_8 _06398_ (.A(_01667_),
    .X(_01668_));
 sky130_fd_sc_hd__and3_2 _06399_ (.A(_01538_),
    .B(_01558_),
    .C(_01573_),
    .X(_01669_));
 sky130_fd_sc_hd__clkbuf_8 _06400_ (.A(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__buf_4 _06401_ (.A(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__and3_2 _06402_ (.A(_01513_),
    .B(_01515_),
    .C(_01553_),
    .X(_01672_));
 sky130_fd_sc_hd__clkbuf_8 _06403_ (.A(_01672_),
    .X(_01673_));
 sky130_fd_sc_hd__clkbuf_8 _06404_ (.A(_01673_),
    .X(_01674_));
 sky130_fd_sc_hd__a22o_1 _06405_ (.A1(\u_rf.reg27_q[0] ),
    .A2(_01671_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[0] ),
    .X(_01675_));
 sky130_fd_sc_hd__a221o_1 _06406_ (.A1(\u_rf.reg0_q[0] ),
    .A2(_01664_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[0] ),
    .C1(_01675_),
    .X(_01676_));
 sky130_fd_sc_hd__or4_1 _06407_ (.A(_01633_),
    .B(_01647_),
    .C(_01661_),
    .D(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__and3b_2 _06408_ (.A_N(_01547_),
    .B(_01517_),
    .C(_01527_),
    .X(_01678_));
 sky130_fd_sc_hd__clkbuf_8 _06409_ (.A(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__buf_4 _06410_ (.A(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__o21a_1 _06411_ (.A1(_01619_),
    .A2(_01677_),
    .B1(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__a221oi_2 _06412_ (.A1(\u_decod.dec0.instr_i[20] ),
    .A2(_01530_),
    .B1(_01550_),
    .B2(\u_decod.rf_ff_res_data_i[0] ),
    .C1(_01681_),
    .Y(_01682_));
 sky130_fd_sc_hd__o21ai_1 _06413_ (.A1(_01511_),
    .A2(_01528_),
    .B1(_01682_),
    .Y(\u_decod.rs2_data_nxt[0] ));
 sky130_fd_sc_hd__and2_1 _06414_ (.A(_01267_),
    .B(_01430_),
    .X(_01683_));
 sky130_fd_sc_hd__inv_2 _06415_ (.A(\u_decod.rs2_data_q[3] ),
    .Y(_01684_));
 sky130_fd_sc_hd__buf_2 _06416_ (.A(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__mux4_1 _06417_ (.A0(_01388_),
    .A1(_01683_),
    .A2(\u_decod.rs1_data_q[8] ),
    .A3(\u_decod.rs1_data_q[24] ),
    .S0(_01446_),
    .S1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _06418_ (.A0(_01471_),
    .A1(_01686_),
    .S(_01464_),
    .X(_01687_));
 sky130_fd_sc_hd__buf_2 _06419_ (.A(_01315_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _06420_ (.A0(_01465_),
    .A1(_01687_),
    .S(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__or2_1 _06421_ (.A(_01474_),
    .B(_01452_),
    .X(_01690_));
 sky130_fd_sc_hd__or2_1 _06422_ (.A(_01493_),
    .B(_01459_),
    .X(_01691_));
 sky130_fd_sc_hd__a21o_1 _06423_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01422_),
    .X(_01692_));
 sky130_fd_sc_hd__o211a_1 _06424_ (.A1(_01479_),
    .A2(_01689_),
    .B1(_01692_),
    .C1(_01441_),
    .X(_01693_));
 sky130_fd_sc_hd__or2_1 _06425_ (.A(_01314_),
    .B(_01316_),
    .X(_01694_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(_01314_),
    .B(_01316_),
    .Y(_01695_));
 sky130_fd_sc_hd__o21a_1 _06427_ (.A1(\u_decod.rs1_data_q[1] ),
    .A2(_01493_),
    .B1(_01431_),
    .X(_01696_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(\u_decod.instr_operation_q[3] ),
    .B(_01259_),
    .Y(_01697_));
 sky130_fd_sc_hd__nor2_1 _06429_ (.A(_01316_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__a32o_1 _06430_ (.A1(\u_decod.rs1_data_q[1] ),
    .A2(_01493_),
    .A3(_01428_),
    .B1(_01484_),
    .B2(\u_decod.pc_q_o[1] ),
    .X(_01699_));
 sky130_fd_sc_hd__or3_1 _06431_ (.A(_01696_),
    .B(_01698_),
    .C(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__a31o_1 _06432_ (.A1(_01694_),
    .A2(_01436_),
    .A3(_01695_),
    .B1(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__clkbuf_4 _06433_ (.A(_01445_),
    .X(_01702_));
 sky130_fd_sc_hd__buf_2 _06434_ (.A(_01494_),
    .X(_01703_));
 sky130_fd_sc_hd__o21a_1 _06435_ (.A1(\u_decod.rs1_data_q[1] ),
    .A2(_01702_),
    .B1(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__o21a_1 _06436_ (.A1(_01455_),
    .A2(_01704_),
    .B1(_01497_),
    .X(_01705_));
 sky130_fd_sc_hd__o21a_1 _06437_ (.A1(_01451_),
    .A2(_01705_),
    .B1(_01500_),
    .X(_01706_));
 sky130_fd_sc_hd__o21a_1 _06438_ (.A1(_01493_),
    .A2(_01706_),
    .B1(_01502_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _06439_ (.A0(_01503_),
    .A1(_01707_),
    .S(_01478_),
    .X(_01708_));
 sky130_fd_sc_hd__a22o_1 _06440_ (.A1(net64),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net50),
    .X(_01709_));
 sky130_fd_sc_hd__a221o_1 _06441_ (.A1(net44),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net41),
    .C1(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__a22o_1 _06442_ (.A1(_01505_),
    .A2(_01708_),
    .B1(_01710_),
    .B2(_01058_),
    .X(_01711_));
 sky130_fd_sc_hd__or3_1 _06443_ (.A(_01693_),
    .B(_01701_),
    .C(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__buf_1 _06444_ (.A(_01712_),
    .X(\u_decod.exe_ff_res_data_i[1] ));
 sky130_fd_sc_hd__nor2_4 _06445_ (.A(_01518_),
    .B(_01527_),
    .Y(_01713_));
 sky130_fd_sc_hd__or2_2 _06446_ (.A(_01206_),
    .B(_01530_),
    .X(_01714_));
 sky130_fd_sc_hd__or2_2 _06447_ (.A(_01205_),
    .B(_01529_),
    .X(_01715_));
 sky130_fd_sc_hd__a22o_1 _06448_ (.A1(\u_decod.dec0.instr_i[8] ),
    .A2(_01226_),
    .B1(_01715_),
    .B2(\u_decod.dec0.instr_i[21] ),
    .X(_01716_));
 sky130_fd_sc_hd__a22o_1 _06449_ (.A1(\u_decod.rf_ff_res_data_i[1] ),
    .A2(_01549_),
    .B1(_01714_),
    .B2(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__a22o_1 _06450_ (.A1(\u_rf.reg16_q[1] ),
    .A2(_01564_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[1] ),
    .X(_01718_));
 sky130_fd_sc_hd__a221o_1 _06451_ (.A1(\u_rf.reg6_q[1] ),
    .A2(_01555_),
    .B1(_01580_),
    .B2(\u_rf.reg30_q[1] ),
    .C1(_01718_),
    .X(_01719_));
 sky130_fd_sc_hd__a22o_1 _06452_ (.A1(\u_rf.reg28_q[1] ),
    .A2(_01624_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[1] ),
    .X(_01720_));
 sky130_fd_sc_hd__a221o_1 _06453_ (.A1(\u_rf.reg1_q[1] ),
    .A2(_01586_),
    .B1(_01615_),
    .B2(\u_rf.reg31_q[1] ),
    .C1(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__a22o_1 _06454_ (.A1(\u_rf.reg10_q[1] ),
    .A2(_01656_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[1] ),
    .X(_01722_));
 sky130_fd_sc_hd__a221o_1 _06455_ (.A1(\u_rf.reg5_q[1] ),
    .A2(_01568_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[1] ),
    .C1(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__a22o_1 _06456_ (.A1(\u_rf.reg13_q[1] ),
    .A2(_01597_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[1] ),
    .X(_01724_));
 sky130_fd_sc_hd__a221o_1 _06457_ (.A1(\u_rf.reg0_q[1] ),
    .A2(_01662_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[1] ),
    .C1(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__or4_1 _06458_ (.A(_01719_),
    .B(_01721_),
    .C(_01723_),
    .D(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__a22o_1 _06459_ (.A1(\u_rf.reg24_q[1] ),
    .A2(_01621_),
    .B1(_01627_),
    .B2(\u_rf.reg29_q[1] ),
    .X(_01727_));
 sky130_fd_sc_hd__a221o_1 _06460_ (.A1(\u_rf.reg25_q[1] ),
    .A2(_01576_),
    .B1(_01630_),
    .B2(\u_rf.reg17_q[1] ),
    .C1(_01727_),
    .X(_01728_));
 sky130_fd_sc_hd__a22o_1 _06461_ (.A1(\u_rf.reg7_q[1] ),
    .A2(_01560_),
    .B1(_01605_),
    .B2(\u_rf.reg3_q[1] ),
    .X(_01729_));
 sky130_fd_sc_hd__a221o_1 _06462_ (.A1(\u_rf.reg19_q[1] ),
    .A2(_01594_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[1] ),
    .C1(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__a22o_1 _06463_ (.A1(\u_rf.reg18_q[1] ),
    .A2(_01591_),
    .B1(_01612_),
    .B2(\u_rf.reg23_q[1] ),
    .X(_01731_));
 sky130_fd_sc_hd__a221o_1 _06464_ (.A1(\u_rf.reg9_q[1] ),
    .A2(_01635_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[1] ),
    .C1(_01731_),
    .X(_01732_));
 sky130_fd_sc_hd__a22o_1 _06465_ (.A1(\u_rf.reg15_q[1] ),
    .A2(_01600_),
    .B1(_01608_),
    .B2(\u_rf.reg12_q[1] ),
    .X(_01733_));
 sky130_fd_sc_hd__a221o_1 _06466_ (.A1(\u_rf.reg11_q[1] ),
    .A2(_01583_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[1] ),
    .C1(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__or4_1 _06467_ (.A(_01728_),
    .B(_01730_),
    .C(_01732_),
    .D(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__o21a_1 _06468_ (.A1(_01726_),
    .A2(_01735_),
    .B1(_01679_),
    .X(_01736_));
 sky130_fd_sc_hd__a211o_1 _06469_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[1] ),
    .B1(_01717_),
    .C1(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__or4_1 _06470_ (.A(_01234_),
    .B(_01079_),
    .C(_01231_),
    .D(_01083_),
    .X(_01738_));
 sky130_fd_sc_hd__o21ai_1 _06471_ (.A1(_01085_),
    .A2(_01738_),
    .B1(_01233_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor4_1 _06472_ (.A(\u_decod.dec0.funct7[3] ),
    .B(\u_decod.dec0.funct7[2] ),
    .C(\u_decod.dec0.funct7[4] ),
    .D(_01081_),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _06473_ (.A(_01197_),
    .B(_01232_),
    .Y(_01741_));
 sky130_fd_sc_hd__and4_1 _06474_ (.A(_01079_),
    .B(_01075_),
    .C(_01740_),
    .D(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__nor4_2 _06475_ (.A(_01089_),
    .B(_01739_),
    .C(_01243_),
    .D(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__inv_2 _06476_ (.A(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _06477_ (.A(\u_decod.rs2_data_nxt[0] ),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__xnor2_1 _06478_ (.A(_01737_),
    .B(_01745_),
    .Y(\u_decod.rs2_data_nxt[1] ));
 sky130_fd_sc_hd__buf_2 _06479_ (.A(_01506_),
    .X(_01746_));
 sky130_fd_sc_hd__buf_2 _06480_ (.A(_01683_),
    .X(_01747_));
 sky130_fd_sc_hd__o21a_1 _06481_ (.A1(_01445_),
    .A2(\u_decod.rs1_data_q[2] ),
    .B1(_01703_),
    .X(_01748_));
 sky130_fd_sc_hd__o21a_1 _06482_ (.A1(_01444_),
    .A2(_01748_),
    .B1(_01497_),
    .X(_01749_));
 sky130_fd_sc_hd__o21a_1 _06483_ (.A1(_01464_),
    .A2(_01749_),
    .B1(_01500_),
    .X(_01750_));
 sky130_fd_sc_hd__mux4_1 _06484_ (.A0(_01747_),
    .A1(_01501_),
    .A2(_01706_),
    .A3(_01750_),
    .S0(_01480_),
    .S1(_01477_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _06485_ (.A0(\u_decod.rs1_data_q[9] ),
    .A1(\u_decod.rs1_data_q[25] ),
    .S(_01702_),
    .X(_01752_));
 sky130_fd_sc_hd__buf_2 _06486_ (.A(_01494_),
    .X(_01753_));
 sky130_fd_sc_hd__o21a_1 _06487_ (.A1(\u_decod.rs1_data_q[17] ),
    .A2(_01446_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _06488_ (.A0(_01752_),
    .A1(_01754_),
    .S(_01467_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(_01453_),
    .A1(_01755_),
    .S(_01464_),
    .X(_01756_));
 sky130_fd_sc_hd__clkbuf_4 _06490_ (.A(_01688_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _06491_ (.A0(_01452_),
    .A1(_01756_),
    .S(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__or2_1 _06492_ (.A(_01424_),
    .B(_01689_),
    .X(_01759_));
 sky130_fd_sc_hd__o211a_1 _06493_ (.A1(_01480_),
    .A2(_01758_),
    .B1(_01759_),
    .C1(_01442_),
    .X(_01760_));
 sky130_fd_sc_hd__a22o_1 _06494_ (.A1(net34),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net51),
    .X(_01761_));
 sky130_fd_sc_hd__a221o_1 _06495_ (.A1(net55),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net42),
    .C1(_01761_),
    .X(_01762_));
 sky130_fd_sc_hd__nand2_4 _06496_ (.A(\u_decod.instr_operation_q[1] ),
    .B(_01259_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand2_4 _06497_ (.A(\u_decod.instr_unit_q[2] ),
    .B(_01056_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_4 _06498_ (.A(\u_decod.instr_operation_q[0] ),
    .B(_01259_),
    .Y(_01765_));
 sky130_fd_sc_hd__and2b_1 _06499_ (.A_N(_01313_),
    .B(_01317_),
    .X(_01766_));
 sky130_fd_sc_hd__a211o_1 _06500_ (.A1(_01318_),
    .A2(_01694_),
    .B1(_01765_),
    .C1(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__o221ai_1 _06501_ (.A1(_01317_),
    .A2(_01763_),
    .B1(_01764_),
    .B2(\u_decod.pc_q_o[2] ),
    .C1(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__a221o_1 _06502_ (.A1(_01317_),
    .A2(_01435_),
    .B1(_01436_),
    .B2(_01319_),
    .C1(_01432_),
    .X(_01769_));
 sky130_fd_sc_hd__and2b_1 _06503_ (.A_N(_01313_),
    .B(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__a211o_1 _06504_ (.A1(_01059_),
    .A2(_01762_),
    .B1(_01768_),
    .C1(_01770_),
    .X(_01771_));
 sky130_fd_sc_hd__a211o_1 _06505_ (.A1(_01746_),
    .A2(_01751_),
    .B1(_01760_),
    .C1(_01771_),
    .X(\u_decod.exe_ff_res_data_i[2] ));
 sky130_fd_sc_hd__clkbuf_4 _06506_ (.A(_01713_),
    .X(_01772_));
 sky130_fd_sc_hd__clkbuf_4 _06507_ (.A(_01714_),
    .X(_01773_));
 sky130_fd_sc_hd__a22o_1 _06508_ (.A1(\u_decod.dec0.instr_i[9] ),
    .A2(_01226_),
    .B1(_01715_),
    .B2(\u_decod.dec0.instr_i[22] ),
    .X(_01774_));
 sky130_fd_sc_hd__a22o_1 _06509_ (.A1(\u_decod.rf_ff_res_data_i[2] ),
    .A2(_01549_),
    .B1(_01773_),
    .B2(_01774_),
    .X(_01775_));
 sky130_fd_sc_hd__clkbuf_8 _06510_ (.A(_01674_),
    .X(_01776_));
 sky130_fd_sc_hd__buf_4 _06511_ (.A(_01616_),
    .X(_01777_));
 sky130_fd_sc_hd__a22o_1 _06512_ (.A1(\u_rf.reg31_q[2] ),
    .A2(_01777_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[2] ),
    .X(_01778_));
 sky130_fd_sc_hd__a221o_1 _06513_ (.A1(\u_rf.reg12_q[2] ),
    .A2(_01610_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[2] ),
    .C1(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__clkbuf_8 _06514_ (.A(_01628_),
    .X(_01780_));
 sky130_fd_sc_hd__a22o_1 _06515_ (.A1(\u_rf.reg14_q[2] ),
    .A2(_01659_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[2] ),
    .X(_01781_));
 sky130_fd_sc_hd__a221o_1 _06516_ (.A1(\u_rf.reg29_q[2] ),
    .A2(_01780_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[2] ),
    .C1(_01781_),
    .X(_01782_));
 sky130_fd_sc_hd__clkbuf_8 _06517_ (.A(_01576_),
    .X(_01783_));
 sky130_fd_sc_hd__clkbuf_8 _06518_ (.A(_01622_),
    .X(_01784_));
 sky130_fd_sc_hd__a22o_1 _06519_ (.A1(\u_rf.reg26_q[2] ),
    .A2(_01642_),
    .B1(_01645_),
    .B2(\u_rf.reg20_q[2] ),
    .X(_01785_));
 sky130_fd_sc_hd__a221o_1 _06520_ (.A1(\u_rf.reg25_q[2] ),
    .A2(_01783_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[2] ),
    .C1(_01785_),
    .X(_01786_));
 sky130_fd_sc_hd__clkbuf_8 _06521_ (.A(_01592_),
    .X(_01787_));
 sky130_fd_sc_hd__a22o_1 _06522_ (.A1(\u_rf.reg30_q[2] ),
    .A2(_01580_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[2] ),
    .X(_01788_));
 sky130_fd_sc_hd__a221o_1 _06523_ (.A1(\u_rf.reg13_q[2] ),
    .A2(_01598_),
    .B1(_01787_),
    .B2(\u_rf.reg18_q[2] ),
    .C1(_01788_),
    .X(_01789_));
 sky130_fd_sc_hd__or3_1 _06524_ (.A(_01782_),
    .B(_01786_),
    .C(_01789_),
    .X(_01790_));
 sky130_fd_sc_hd__clkbuf_8 _06525_ (.A(_01656_),
    .X(_01791_));
 sky130_fd_sc_hd__a22o_1 _06526_ (.A1(\u_rf.reg6_q[2] ),
    .A2(_01556_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[2] ),
    .X(_01792_));
 sky130_fd_sc_hd__a221o_1 _06527_ (.A1(\u_rf.reg23_q[2] ),
    .A2(_01613_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[2] ),
    .C1(_01792_),
    .X(_01793_));
 sky130_fd_sc_hd__a22o_1 _06528_ (.A1(\u_rf.reg1_q[2] ),
    .A2(_01586_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[2] ),
    .X(_01794_));
 sky130_fd_sc_hd__a221o_1 _06529_ (.A1(\u_rf.reg11_q[2] ),
    .A2(_01584_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[2] ),
    .C1(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__a22o_1 _06530_ (.A1(\u_rf.reg7_q[2] ),
    .A2(_01561_),
    .B1(_01606_),
    .B2(\u_rf.reg3_q[2] ),
    .X(_01796_));
 sky130_fd_sc_hd__a221o_1 _06531_ (.A1(\u_rf.reg0_q[2] ),
    .A2(_01663_),
    .B1(_01601_),
    .B2(\u_rf.reg15_q[2] ),
    .C1(_01796_),
    .X(_01797_));
 sky130_fd_sc_hd__a22o_1 _06532_ (.A1(\u_rf.reg16_q[2] ),
    .A2(_01565_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[2] ),
    .X(_01798_));
 sky130_fd_sc_hd__a221o_1 _06533_ (.A1(\u_rf.reg5_q[2] ),
    .A2(_01569_),
    .B1(_01595_),
    .B2(\u_rf.reg19_q[2] ),
    .C1(_01798_),
    .X(_01799_));
 sky130_fd_sc_hd__or4_1 _06534_ (.A(_01793_),
    .B(_01795_),
    .C(_01797_),
    .D(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__o31a_1 _06535_ (.A1(_01779_),
    .A2(_01790_),
    .A3(_01800_),
    .B1(_01680_),
    .X(_01801_));
 sky130_fd_sc_hd__a211o_1 _06536_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[2] ),
    .B1(_01775_),
    .C1(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__inv_2 _06537_ (.A(_01737_),
    .Y(_01803_));
 sky130_fd_sc_hd__o211a_1 _06538_ (.A1(_01511_),
    .A2(_01528_),
    .B1(_01682_),
    .C1(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__nor2_1 _06539_ (.A(net201),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__xor2_1 _06540_ (.A(_01802_),
    .B(_01805_),
    .X(\u_decod.rs2_data_nxt[2] ));
 sky130_fd_sc_hd__mux4_1 _06541_ (.A0(_01384_),
    .A1(_01683_),
    .A2(_01302_),
    .A3(\u_decod.rs1_data_q[26] ),
    .S0(_01446_),
    .S1(_01685_),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _06542_ (.A0(_01463_),
    .A1(_01806_),
    .S(_01451_),
    .X(_01807_));
 sky130_fd_sc_hd__mux2_1 _06543_ (.A0(_01687_),
    .A1(_01807_),
    .S(_01688_),
    .X(_01808_));
 sky130_fd_sc_hd__or2_1 _06544_ (.A(_01479_),
    .B(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__o211a_1 _06545_ (.A1(_01424_),
    .A2(_01758_),
    .B1(_01809_),
    .C1(_01441_),
    .X(_01810_));
 sky130_fd_sc_hd__nor2_1 _06546_ (.A(_01313_),
    .B(_01319_),
    .Y(_01811_));
 sky130_fd_sc_hd__and2_1 _06547_ (.A(\u_decod.rs1_data_q[3] ),
    .B(_01468_),
    .X(_01812_));
 sky130_fd_sc_hd__nor2_1 _06548_ (.A(_01812_),
    .B(_01312_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21oi_1 _06549_ (.A1(_01811_),
    .A2(_01813_),
    .B1(_01765_),
    .Y(_01814_));
 sky130_fd_sc_hd__o21a_1 _06550_ (.A1(_01811_),
    .A2(_01813_),
    .B1(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__nand2_1 _06551_ (.A(\u_decod.pc_q_o[2] ),
    .B(\u_decod.pc_q_o[3] ),
    .Y(_01816_));
 sky130_fd_sc_hd__or2_1 _06552_ (.A(\u_decod.pc_q_o[2] ),
    .B(\u_decod.pc_q_o[3] ),
    .X(_01817_));
 sky130_fd_sc_hd__a32o_1 _06553_ (.A1(_01484_),
    .A2(_01816_),
    .A3(_01817_),
    .B1(_01813_),
    .B2(_01435_),
    .X(_01818_));
 sky130_fd_sc_hd__nand2_2 _06554_ (.A(_01430_),
    .B(_01259_),
    .Y(_01819_));
 sky130_fd_sc_hd__clkbuf_4 _06555_ (.A(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__o22a_1 _06556_ (.A1(_01320_),
    .A2(_01763_),
    .B1(_01820_),
    .B2(_01312_),
    .X(_01821_));
 sky130_fd_sc_hd__or3b_1 _06557_ (.A(_01815_),
    .B(_01818_),
    .C_N(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__o21a_1 _06558_ (.A1(_01702_),
    .A2(\u_decod.rs1_data_q[3] ),
    .B1(_01703_),
    .X(_01823_));
 sky130_fd_sc_hd__o21a_1 _06559_ (.A1(_01444_),
    .A2(_01823_),
    .B1(_01497_),
    .X(_01824_));
 sky130_fd_sc_hd__o21a_1 _06560_ (.A1(_01464_),
    .A2(_01824_),
    .B1(_01500_),
    .X(_01825_));
 sky130_fd_sc_hd__mux4_1 _06561_ (.A0(_01501_),
    .A1(_01706_),
    .A2(_01750_),
    .A3(_01825_),
    .S0(_01479_),
    .S1(_01476_),
    .X(_01826_));
 sky130_fd_sc_hd__a22o_1 _06562_ (.A1(net35),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net52),
    .X(_01827_));
 sky130_fd_sc_hd__a221o_1 _06563_ (.A1(net58),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net43),
    .C1(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__a22o_1 _06564_ (.A1(_01506_),
    .A2(_01826_),
    .B1(_01828_),
    .B2(_01059_),
    .X(_01829_));
 sky130_fd_sc_hd__or3_1 _06565_ (.A(_01810_),
    .B(_01822_),
    .C(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__buf_1 _06566_ (.A(_01830_),
    .X(\u_decod.exe_ff_res_data_i[3] ));
 sky130_fd_sc_hd__a22o_1 _06567_ (.A1(\u_decod.dec0.instr_i[10] ),
    .A2(_01226_),
    .B1(_01715_),
    .B2(\u_decod.dec0.instr_i[23] ),
    .X(_01831_));
 sky130_fd_sc_hd__a22o_1 _06568_ (.A1(\u_decod.rf_ff_res_data_i[3] ),
    .A2(_01549_),
    .B1(_01773_),
    .B2(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__a22o_1 _06569_ (.A1(\u_rf.reg25_q[3] ),
    .A2(_01575_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[3] ),
    .X(_01833_));
 sky130_fd_sc_hd__a221o_1 _06570_ (.A1(\u_rf.reg16_q[3] ),
    .A2(_01564_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[3] ),
    .C1(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__a22o_1 _06571_ (.A1(\u_rf.reg12_q[3] ),
    .A2(_01608_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[3] ),
    .X(_01835_));
 sky130_fd_sc_hd__a221o_1 _06572_ (.A1(\u_rf.reg3_q[3] ),
    .A2(_01605_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[3] ),
    .C1(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__a22o_1 _06573_ (.A1(\u_rf.reg6_q[3] ),
    .A2(_01555_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[3] ),
    .X(_01837_));
 sky130_fd_sc_hd__a221o_1 _06574_ (.A1(\u_rf.reg29_q[3] ),
    .A2(_01628_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[3] ),
    .C1(_01837_),
    .X(_01838_));
 sky130_fd_sc_hd__a22o_1 _06575_ (.A1(\u_rf.reg15_q[3] ),
    .A2(_01600_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[3] ),
    .X(_01839_));
 sky130_fd_sc_hd__a221o_1 _06576_ (.A1(\u_rf.reg5_q[3] ),
    .A2(_01569_),
    .B1(_01561_),
    .B2(\u_rf.reg7_q[3] ),
    .C1(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__or4_1 _06577_ (.A(_01834_),
    .B(_01836_),
    .C(_01838_),
    .D(_01840_),
    .X(_01841_));
 sky130_fd_sc_hd__a22o_1 _06578_ (.A1(\u_rf.reg19_q[3] ),
    .A2(_01594_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[3] ),
    .X(_01842_));
 sky130_fd_sc_hd__a221o_1 _06579_ (.A1(\u_rf.reg11_q[3] ),
    .A2(_01583_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[3] ),
    .C1(_01842_),
    .X(_01843_));
 sky130_fd_sc_hd__a22o_1 _06580_ (.A1(\u_rf.reg31_q[3] ),
    .A2(_01615_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[3] ),
    .X(_01844_));
 sky130_fd_sc_hd__a221o_1 _06581_ (.A1(\u_rf.reg23_q[3] ),
    .A2(_01613_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[3] ),
    .C1(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__a22o_1 _06582_ (.A1(\u_rf.reg30_q[3] ),
    .A2(_01579_),
    .B1(_01597_),
    .B2(\u_rf.reg13_q[3] ),
    .X(_01846_));
 sky130_fd_sc_hd__a221o_1 _06583_ (.A1(\u_rf.reg0_q[3] ),
    .A2(_01663_),
    .B1(_01645_),
    .B2(\u_rf.reg20_q[3] ),
    .C1(_01846_),
    .X(_01847_));
 sky130_fd_sc_hd__a22o_1 _06584_ (.A1(\u_rf.reg9_q[3] ),
    .A2(_01635_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[3] ),
    .X(_01848_));
 sky130_fd_sc_hd__a221o_1 _06585_ (.A1(\u_rf.reg1_q[3] ),
    .A2(_01587_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[3] ),
    .C1(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__or4_1 _06586_ (.A(_01843_),
    .B(_01845_),
    .C(_01847_),
    .D(_01849_),
    .X(_01850_));
 sky130_fd_sc_hd__or2_1 _06587_ (.A(_01841_),
    .B(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__and2_1 _06588_ (.A(_01680_),
    .B(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__a211o_1 _06589_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[3] ),
    .B1(_01832_),
    .C1(_01852_),
    .X(_01853_));
 sky130_fd_sc_hd__o21ai_1 _06590_ (.A1(_01802_),
    .A2(_01805_),
    .B1(_01744_),
    .Y(_01854_));
 sky130_fd_sc_hd__xnor2_1 _06591_ (.A(_01853_),
    .B(_01854_),
    .Y(\u_decod.rs2_data_nxt[3] ));
 sky130_fd_sc_hd__a22o_1 _06592_ (.A1(net36),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net53),
    .X(_01855_));
 sky130_fd_sc_hd__a221o_1 _06593_ (.A1(net59),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net45),
    .C1(_01855_),
    .X(_01856_));
 sky130_fd_sc_hd__a21oi_1 _06594_ (.A1(\u_decod.pc_q_o[2] ),
    .A2(\u_decod.pc_q_o[3] ),
    .B1(\u_decod.pc_q_o[4] ),
    .Y(_01857_));
 sky130_fd_sc_hd__a31o_1 _06595_ (.A1(\u_decod.pc_q_o[2] ),
    .A2(\u_decod.pc_q_o[3] ),
    .A3(\u_decod.pc_q_o[4] ),
    .B1(_01764_),
    .X(_01858_));
 sky130_fd_sc_hd__o22ai_1 _06596_ (.A1(_01323_),
    .A2(_01763_),
    .B1(_01857_),
    .B2(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _06597_ (.A(_01321_),
    .B(_01324_),
    .Y(_01860_));
 sky130_fd_sc_hd__or2_1 _06598_ (.A(_01321_),
    .B(_01324_),
    .X(_01861_));
 sky130_fd_sc_hd__a32o_1 _06599_ (.A1(_01860_),
    .A2(_01436_),
    .A3(_01861_),
    .B1(_01435_),
    .B2(_01324_),
    .X(_01862_));
 sky130_fd_sc_hd__a211o_1 _06600_ (.A1(_01322_),
    .A2(_01432_),
    .B1(_01859_),
    .C1(_01862_),
    .X(_01863_));
 sky130_fd_sc_hd__and2_1 _06601_ (.A(_01322_),
    .B(_01494_),
    .X(_01864_));
 sky130_fd_sc_hd__o21a_1 _06602_ (.A1(\u_decod.rs2_data_q[3] ),
    .A2(_01864_),
    .B1(_01497_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _06603_ (.A0(_01499_),
    .A1(_01865_),
    .S(_01458_),
    .X(_01866_));
 sky130_fd_sc_hd__mux4_1 _06604_ (.A0(_01706_),
    .A1(_01750_),
    .A2(_01825_),
    .A3(_01866_),
    .S0(_01479_),
    .S1(_01476_),
    .X(_01867_));
 sky130_fd_sc_hd__mux4_1 _06605_ (.A0(\u_decod.rs1_data_q[19] ),
    .A1(_01683_),
    .A2(\u_decod.rs1_data_q[11] ),
    .A3(\u_decod.rs1_data_q[27] ),
    .S0(_01702_),
    .S1(_01684_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _06606_ (.A0(_01449_),
    .A1(_01868_),
    .S(_01464_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _06607_ (.A0(_01756_),
    .A1(_01869_),
    .S(_01688_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _06608_ (.A0(_01808_),
    .A1(_01870_),
    .S(_01423_),
    .X(_01871_));
 sky130_fd_sc_hd__a22o_1 _06609_ (.A1(_01506_),
    .A2(_01867_),
    .B1(_01871_),
    .B2(_01442_),
    .X(_01872_));
 sky130_fd_sc_hd__a211oi_2 _06610_ (.A1(net133),
    .A2(_01856_),
    .B1(_01863_),
    .C1(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__inv_2 _06611_ (.A(_01873_),
    .Y(\u_decod.exe_ff_res_data_i[4] ));
 sky130_fd_sc_hd__a22o_1 _06612_ (.A1(\u_decod.dec0.instr_i[11] ),
    .A2(_01226_),
    .B1(_01715_),
    .B2(_01572_),
    .X(_01874_));
 sky130_fd_sc_hd__a22o_1 _06613_ (.A1(\u_rf.reg26_q[4] ),
    .A2(_01641_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[4] ),
    .X(_01875_));
 sky130_fd_sc_hd__a221o_1 _06614_ (.A1(\u_rf.reg25_q[4] ),
    .A2(_01575_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[4] ),
    .C1(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__a22o_1 _06615_ (.A1(\u_rf.reg30_q[4] ),
    .A2(_01579_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[4] ),
    .X(_01877_));
 sky130_fd_sc_hd__a221o_1 _06616_ (.A1(\u_rf.reg13_q[4] ),
    .A2(_01597_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[4] ),
    .C1(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__a22o_1 _06617_ (.A1(\u_rf.reg31_q[4] ),
    .A2(_01615_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[4] ),
    .X(_01879_));
 sky130_fd_sc_hd__a221o_1 _06618_ (.A1(\u_rf.reg12_q[4] ),
    .A2(_01608_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[4] ),
    .C1(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__a22o_1 _06619_ (.A1(\u_rf.reg14_q[4] ),
    .A2(_01658_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[4] ),
    .X(_01881_));
 sky130_fd_sc_hd__a221o_1 _06620_ (.A1(\u_rf.reg29_q[4] ),
    .A2(_01628_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[4] ),
    .C1(_01881_),
    .X(_01882_));
 sky130_fd_sc_hd__or4_1 _06621_ (.A(_01876_),
    .B(_01878_),
    .C(_01880_),
    .D(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__a22o_1 _06622_ (.A1(\u_rf.reg6_q[4] ),
    .A2(_01555_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[4] ),
    .X(_01884_));
 sky130_fd_sc_hd__a221o_1 _06623_ (.A1(\u_rf.reg23_q[4] ),
    .A2(_01613_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[4] ),
    .C1(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__a22o_1 _06624_ (.A1(\u_rf.reg1_q[4] ),
    .A2(_01586_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[4] ),
    .X(_01886_));
 sky130_fd_sc_hd__a221o_1 _06625_ (.A1(\u_rf.reg11_q[4] ),
    .A2(_01583_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[4] ),
    .C1(_01886_),
    .X(_01887_));
 sky130_fd_sc_hd__a22o_1 _06626_ (.A1(\u_rf.reg7_q[4] ),
    .A2(_01560_),
    .B1(_01605_),
    .B2(\u_rf.reg3_q[4] ),
    .X(_01888_));
 sky130_fd_sc_hd__a221o_1 _06627_ (.A1(\u_rf.reg0_q[4] ),
    .A2(_01662_),
    .B1(_01601_),
    .B2(\u_rf.reg15_q[4] ),
    .C1(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__a22o_1 _06628_ (.A1(\u_rf.reg16_q[4] ),
    .A2(_01564_),
    .B1(_01630_),
    .B2(\u_rf.reg17_q[4] ),
    .X(_01890_));
 sky130_fd_sc_hd__a221o_1 _06629_ (.A1(\u_rf.reg5_q[4] ),
    .A2(_01569_),
    .B1(_01594_),
    .B2(\u_rf.reg19_q[4] ),
    .C1(_01890_),
    .X(_01891_));
 sky130_fd_sc_hd__or4_1 _06630_ (.A(_01885_),
    .B(_01887_),
    .C(_01889_),
    .D(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__o21a_1 _06631_ (.A1(_01883_),
    .A2(_01892_),
    .B1(_01679_),
    .X(_01893_));
 sky130_fd_sc_hd__a221o_1 _06632_ (.A1(\u_decod.rf_ff_res_data_i[4] ),
    .A2(_01549_),
    .B1(_01714_),
    .B2(_01874_),
    .C1(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__a21o_1 _06633_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[4] ),
    .B1(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__and3_1 _06634_ (.A(_01075_),
    .B(_01740_),
    .C(_01741_),
    .X(_01896_));
 sky130_fd_sc_hd__a221o_4 _06635_ (.A1(_01093_),
    .A2(_01090_),
    .B1(_01896_),
    .B2(_01079_),
    .C1(_01237_),
    .X(_01897_));
 sky130_fd_sc_hd__nor2_1 _06636_ (.A(_01802_),
    .B(_01853_),
    .Y(_01898_));
 sky130_fd_sc_hd__nand2_1 _06637_ (.A(_01804_),
    .B(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__nand2_1 _06638_ (.A(_01897_),
    .B(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__xnor2_1 _06639_ (.A(_01895_),
    .B(_01900_),
    .Y(\u_decod.rs2_data_nxt[4] ));
 sky130_fd_sc_hd__a21oi_1 _06640_ (.A1(_01323_),
    .A2(_01860_),
    .B1(_01311_),
    .Y(_01901_));
 sky130_fd_sc_hd__a31o_1 _06641_ (.A1(_01311_),
    .A2(_01323_),
    .A3(_01860_),
    .B1(_01765_),
    .X(_01902_));
 sky130_fd_sc_hd__o21a_1 _06642_ (.A1(\u_decod.rs1_data_q[5] ),
    .A2(_01702_),
    .B1(_01703_),
    .X(_01903_));
 sky130_fd_sc_hd__o21a_1 _06643_ (.A1(_01444_),
    .A2(_01903_),
    .B1(_01497_),
    .X(_01904_));
 sky130_fd_sc_hd__clkbuf_4 _06644_ (.A(_01458_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _06645_ (.A0(_01705_),
    .A1(_01904_),
    .S(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__mux4_1 _06646_ (.A0(_01750_),
    .A1(_01825_),
    .A2(_01866_),
    .A3(_01906_),
    .S0(_01478_),
    .S1(_01475_),
    .X(_01907_));
 sky130_fd_sc_hd__nand2_1 _06647_ (.A(_01505_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__mux4_1 _06648_ (.A0(_01363_),
    .A1(_01683_),
    .A2(_01297_),
    .A3(\u_decod.rs1_data_q[28] ),
    .S0(_01446_),
    .S1(_01685_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _06649_ (.A0(_01686_),
    .A1(_01909_),
    .S(_01450_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _06650_ (.A0(_01807_),
    .A1(_01910_),
    .S(_01688_),
    .X(_01911_));
 sky130_fd_sc_hd__o21a_1 _06651_ (.A1(_01479_),
    .A2(_01911_),
    .B1(_01441_),
    .X(_01912_));
 sky130_fd_sc_hd__o21ai_1 _06652_ (.A1(_01423_),
    .A2(_01870_),
    .B1(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__a22o_1 _06653_ (.A1(net37),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net54),
    .X(_01914_));
 sky130_fd_sc_hd__a221o_1 _06654_ (.A1(net60),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net46),
    .C1(_01914_),
    .X(_01915_));
 sky130_fd_sc_hd__nand2_1 _06655_ (.A(_01058_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__and4_1 _06656_ (.A(\u_decod.pc_q_o[2] ),
    .B(\u_decod.pc_q_o[3] ),
    .C(\u_decod.pc_q_o[4] ),
    .D(\u_decod.pc_q_o[5] ),
    .X(_01917_));
 sky130_fd_sc_hd__a31o_1 _06657_ (.A1(\u_decod.pc_q_o[2] ),
    .A2(\u_decod.pc_q_o[3] ),
    .A3(\u_decod.pc_q_o[4] ),
    .B1(\u_decod.pc_q_o[5] ),
    .X(_01918_));
 sky130_fd_sc_hd__or3b_1 _06658_ (.A(_01764_),
    .B(_01917_),
    .C_N(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__o22a_1 _06659_ (.A1(_01309_),
    .A2(_01819_),
    .B1(_01697_),
    .B2(_01311_),
    .X(_01920_));
 sky130_fd_sc_hd__o2111a_1 _06660_ (.A1(_01310_),
    .A2(_01763_),
    .B1(_01916_),
    .C1(_01919_),
    .D1(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__and3_1 _06661_ (.A(_01908_),
    .B(_01913_),
    .C(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__o21a_1 _06662_ (.A1(_01901_),
    .A2(_01902_),
    .B1(_01922_),
    .X(_01923_));
 sky130_fd_sc_hd__inv_2 _06663_ (.A(_01923_),
    .Y(\u_decod.exe_ff_res_data_i[5] ));
 sky130_fd_sc_hd__a22o_1 _06664_ (.A1(\u_rf.reg30_q[5] ),
    .A2(_01578_),
    .B1(_01599_),
    .B2(\u_rf.reg15_q[5] ),
    .X(_01924_));
 sky130_fd_sc_hd__a221o_1 _06665_ (.A1(\u_rf.reg24_q[5] ),
    .A2(_01621_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[5] ),
    .C1(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__a22o_1 _06666_ (.A1(\u_rf.reg28_q[5] ),
    .A2(_01624_),
    .B1(_01665_),
    .B2(\u_rf.reg8_q[5] ),
    .X(_01926_));
 sky130_fd_sc_hd__a221o_1 _06667_ (.A1(\u_rf.reg25_q[5] ),
    .A2(_01575_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[5] ),
    .C1(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__a22o_1 _06668_ (.A1(\u_rf.reg19_q[5] ),
    .A2(_01593_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[5] ),
    .X(_01928_));
 sky130_fd_sc_hd__a221o_1 _06669_ (.A1(\u_rf.reg26_q[5] ),
    .A2(_01641_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[5] ),
    .C1(_01928_),
    .X(_01929_));
 sky130_fd_sc_hd__a22o_1 _06670_ (.A1(\u_rf.reg1_q[5] ),
    .A2(_01586_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[5] ),
    .X(_01930_));
 sky130_fd_sc_hd__a221o_1 _06671_ (.A1(\u_rf.reg18_q[5] ),
    .A2(_01591_),
    .B1(_01612_),
    .B2(\u_rf.reg23_q[5] ),
    .C1(_01930_),
    .X(_01931_));
 sky130_fd_sc_hd__or4_1 _06672_ (.A(_01925_),
    .B(_01927_),
    .C(_01929_),
    .D(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__a22o_1 _06673_ (.A1(\u_rf.reg12_q[5] ),
    .A2(_01607_),
    .B1(_01637_),
    .B2(\u_rf.reg21_q[5] ),
    .X(_01933_));
 sky130_fd_sc_hd__a221o_1 _06674_ (.A1(\u_rf.reg16_q[5] ),
    .A2(_01564_),
    .B1(_01615_),
    .B2(\u_rf.reg31_q[5] ),
    .C1(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__a22o_1 _06675_ (.A1(\u_rf.reg13_q[5] ),
    .A2(_01596_),
    .B1(_01626_),
    .B2(\u_rf.reg29_q[5] ),
    .X(_01935_));
 sky130_fd_sc_hd__a221o_1 _06676_ (.A1(\u_rf.reg17_q[5] ),
    .A2(_01630_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[5] ),
    .C1(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__a22o_1 _06677_ (.A1(\u_rf.reg7_q[5] ),
    .A2(_01560_),
    .B1(_01604_),
    .B2(\u_rf.reg3_q[5] ),
    .X(_01937_));
 sky130_fd_sc_hd__a221o_1 _06678_ (.A1(\u_rf.reg6_q[5] ),
    .A2(_01555_),
    .B1(_01583_),
    .B2(\u_rf.reg11_q[5] ),
    .C1(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__a22o_1 _06679_ (.A1(\u_rf.reg0_q[5] ),
    .A2(_01662_),
    .B1(_01568_),
    .B2(\u_rf.reg5_q[5] ),
    .X(_01939_));
 sky130_fd_sc_hd__a221o_1 _06680_ (.A1(\u_rf.reg10_q[5] ),
    .A2(_01656_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[5] ),
    .C1(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__or4_1 _06681_ (.A(_01934_),
    .B(_01936_),
    .C(_01938_),
    .D(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__o21a_1 _06682_ (.A1(_01932_),
    .A2(_01941_),
    .B1(_01678_),
    .X(_01942_));
 sky130_fd_sc_hd__a221o_1 _06683_ (.A1(\u_decod.dec0.funct7[0] ),
    .A2(_01530_),
    .B1(_01549_),
    .B2(\u_decod.rf_ff_res_data_i[5] ),
    .C1(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__a21o_1 _06684_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[5] ),
    .B1(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__nor2_1 _06685_ (.A(_01895_),
    .B(_01899_),
    .Y(_01945_));
 sky130_fd_sc_hd__or2_1 _06686_ (.A(_01743_),
    .B(_01945_),
    .X(_01946_));
 sky130_fd_sc_hd__xnor2_1 _06687_ (.A(_01944_),
    .B(_01946_),
    .Y(\u_decod.rs2_data_nxt[5] ));
 sky130_fd_sc_hd__o21a_1 _06688_ (.A1(_01311_),
    .A2(_01860_),
    .B1(_01333_),
    .X(_01947_));
 sky130_fd_sc_hd__xor2_1 _06689_ (.A(_01330_),
    .B(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _06690_ (.A0(\u_decod.rs1_data_q[13] ),
    .A1(\u_decod.rs1_data_q[29] ),
    .S(_01702_),
    .X(_01949_));
 sky130_fd_sc_hd__o21a_1 _06691_ (.A1(\u_decod.rs1_data_q[21] ),
    .A2(_01446_),
    .B1(_01753_),
    .X(_01950_));
 sky130_fd_sc_hd__mux4_1 _06692_ (.A0(_01949_),
    .A1(_01752_),
    .A2(_01950_),
    .A3(_01754_),
    .S0(_01457_),
    .S1(_01460_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _06693_ (.A0(_01869_),
    .A1(_01951_),
    .S(_01688_),
    .X(_01952_));
 sky130_fd_sc_hd__mux2_1 _06694_ (.A0(_01911_),
    .A1(_01952_),
    .S(_01423_),
    .X(_01953_));
 sky130_fd_sc_hd__nand2_1 _06695_ (.A(_01442_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__o21a_1 _06696_ (.A1(\u_decod.rs1_data_q[6] ),
    .A2(_01445_),
    .B1(_01703_),
    .X(_01955_));
 sky130_fd_sc_hd__o211a_1 _06697_ (.A1(\u_decod.rs2_data_q[3] ),
    .A2(_01955_),
    .B1(_01497_),
    .C1(_01457_),
    .X(_01956_));
 sky130_fd_sc_hd__a21o_1 _06698_ (.A1(_01450_),
    .A2(_01749_),
    .B1(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__mux4_1 _06699_ (.A0(_01825_),
    .A1(_01866_),
    .A2(_01906_),
    .A3(_01957_),
    .S0(_01479_),
    .S1(_01476_),
    .X(_01958_));
 sky130_fd_sc_hd__a22o_1 _06700_ (.A1(net38),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net56),
    .X(_01959_));
 sky130_fd_sc_hd__a221o_1 _06701_ (.A1(net61),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net47),
    .C1(_01959_),
    .X(_01960_));
 sky130_fd_sc_hd__or2_1 _06702_ (.A(\u_decod.rs2_data_q[6] ),
    .B(\u_decod.rs1_data_q[6] ),
    .X(_01961_));
 sky130_fd_sc_hd__or2_1 _06703_ (.A(\u_decod.pc_q_o[6] ),
    .B(_01917_),
    .X(_01962_));
 sky130_fd_sc_hd__nand2_1 _06704_ (.A(\u_decod.pc_q_o[6] ),
    .B(_01917_),
    .Y(_01963_));
 sky130_fd_sc_hd__a32o_1 _06705_ (.A1(_01484_),
    .A2(_01962_),
    .A3(_01963_),
    .B1(_01428_),
    .B2(_01329_),
    .X(_01964_));
 sky130_fd_sc_hd__a221o_1 _06706_ (.A1(_01961_),
    .A2(_01431_),
    .B1(_01434_),
    .B2(_01330_),
    .C1(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__a21o_1 _06707_ (.A1(_01058_),
    .A2(_01960_),
    .B1(_01965_),
    .X(_01966_));
 sky130_fd_sc_hd__a21oi_1 _06708_ (.A1(_01506_),
    .A2(_01958_),
    .B1(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__o211a_1 _06709_ (.A1(_01765_),
    .A2(_01948_),
    .B1(_01954_),
    .C1(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__inv_2 _06710_ (.A(_01968_),
    .Y(\u_decod.exe_ff_res_data_i[6] ));
 sky130_fd_sc_hd__a22o_1 _06711_ (.A1(\u_rf.reg9_q[6] ),
    .A2(_01635_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[6] ),
    .X(_01969_));
 sky130_fd_sc_hd__a221o_1 _06712_ (.A1(\u_rf.reg11_q[6] ),
    .A2(_01583_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[6] ),
    .C1(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__a22o_1 _06713_ (.A1(\u_rf.reg17_q[6] ),
    .A2(_01629_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[6] ),
    .X(_01971_));
 sky130_fd_sc_hd__a221o_1 _06714_ (.A1(\u_rf.reg3_q[6] ),
    .A2(_01605_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[6] ),
    .C1(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__a22o_1 _06715_ (.A1(\u_rf.reg18_q[6] ),
    .A2(_01591_),
    .B1(_01669_),
    .B2(\u_rf.reg27_q[6] ),
    .X(_01973_));
 sky130_fd_sc_hd__a221o_1 _06716_ (.A1(\u_rf.reg7_q[6] ),
    .A2(_01560_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[6] ),
    .C1(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__a22o_1 _06717_ (.A1(\u_rf.reg23_q[6] ),
    .A2(_01611_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[6] ),
    .X(_01975_));
 sky130_fd_sc_hd__a221o_1 _06718_ (.A1(\u_rf.reg16_q[6] ),
    .A2(_01564_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[6] ),
    .C1(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__or4_1 _06719_ (.A(_01970_),
    .B(_01972_),
    .C(_01974_),
    .D(_01976_),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_1 _06720_ (.A1(\u_rf.reg1_q[6] ),
    .A2(_01586_),
    .B1(_01575_),
    .B2(\u_rf.reg25_q[6] ),
    .X(_01978_));
 sky130_fd_sc_hd__a221o_1 _06721_ (.A1(\u_rf.reg13_q[6] ),
    .A2(_01597_),
    .B1(_01600_),
    .B2(\u_rf.reg15_q[6] ),
    .C1(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__a22o_1 _06722_ (.A1(\u_rf.reg19_q[6] ),
    .A2(_01593_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[6] ),
    .X(_01980_));
 sky130_fd_sc_hd__a221o_1 _06723_ (.A1(\u_rf.reg0_q[6] ),
    .A2(_01662_),
    .B1(_01627_),
    .B2(\u_rf.reg29_q[6] ),
    .C1(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__a22o_1 _06724_ (.A1(\u_rf.reg31_q[6] ),
    .A2(_01615_),
    .B1(_01648_),
    .B2(\u_rf.reg4_q[6] ),
    .X(_01982_));
 sky130_fd_sc_hd__a221o_1 _06725_ (.A1(\u_rf.reg5_q[6] ),
    .A2(_01568_),
    .B1(_01555_),
    .B2(\u_rf.reg6_q[6] ),
    .C1(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__a22o_1 _06726_ (.A1(\u_rf.reg24_q[6] ),
    .A2(_01621_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[6] ),
    .X(_01984_));
 sky130_fd_sc_hd__a221o_1 _06727_ (.A1(\u_rf.reg30_q[6] ),
    .A2(_01579_),
    .B1(_01608_),
    .B2(\u_rf.reg12_q[6] ),
    .C1(_01984_),
    .X(_01985_));
 sky130_fd_sc_hd__or4_1 _06728_ (.A(_01979_),
    .B(_01981_),
    .C(_01983_),
    .D(_01985_),
    .X(_01986_));
 sky130_fd_sc_hd__or2_1 _06729_ (.A(_01977_),
    .B(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__a22o_1 _06730_ (.A1(\u_decod.dec0.funct7[1] ),
    .A2(_01530_),
    .B1(_01548_),
    .B2(\u_decod.rf_ff_res_data_i[6] ),
    .X(_01988_));
 sky130_fd_sc_hd__a21o_1 _06731_ (.A1(_01679_),
    .A2(_01987_),
    .B1(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__a21o_1 _06732_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[6] ),
    .B1(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__a21boi_1 _06733_ (.A1(_01744_),
    .A2(_01944_),
    .B1_N(_01946_),
    .Y(_01991_));
 sky130_fd_sc_hd__xnor2_1 _06734_ (.A(_01990_),
    .B(_01991_),
    .Y(\u_decod.rs2_data_nxt[6] ));
 sky130_fd_sc_hd__o21ba_1 _06735_ (.A1(_01328_),
    .A2(_01947_),
    .B1_N(_01329_),
    .X(_01992_));
 sky130_fd_sc_hd__xor2_1 _06736_ (.A(_01327_),
    .B(_01992_),
    .X(_01993_));
 sky130_fd_sc_hd__mux4_1 _06737_ (.A0(\u_decod.rs1_data_q[22] ),
    .A1(_01683_),
    .A2(_01292_),
    .A3(\u_decod.rs1_data_q[30] ),
    .S0(_01446_),
    .S1(_01684_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _06738_ (.A0(_01806_),
    .A1(_01994_),
    .S(_01450_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _06739_ (.A0(_01910_),
    .A1(_01995_),
    .S(_01315_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _06740_ (.A0(_01952_),
    .A1(_01996_),
    .S(_01423_),
    .X(_01997_));
 sky130_fd_sc_hd__nand2_1 _06741_ (.A(_01442_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__mux2_1 _06742_ (.A0(_01866_),
    .A1(_01957_),
    .S(_01476_),
    .X(_01999_));
 sky130_fd_sc_hd__o21a_1 _06743_ (.A1(\u_decod.rs1_data_q[7] ),
    .A2(_01702_),
    .B1(_01703_),
    .X(_02000_));
 sky130_fd_sc_hd__o21a_1 _06744_ (.A1(_01444_),
    .A2(_02000_),
    .B1(_01497_),
    .X(_02001_));
 sky130_fd_sc_hd__mux4_1 _06745_ (.A0(_01705_),
    .A1(_01824_),
    .A2(_01904_),
    .A3(_02001_),
    .S0(_01474_),
    .S1(_01457_),
    .X(_02002_));
 sky130_fd_sc_hd__o21a_1 _06746_ (.A1(_01424_),
    .A2(_02002_),
    .B1(_01506_),
    .X(_02003_));
 sky130_fd_sc_hd__o21ai_1 _06747_ (.A1(_01480_),
    .A2(_01999_),
    .B1(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a21oi_1 _06748_ (.A1(\u_decod.pc_q_o[6] ),
    .A2(_01917_),
    .B1(\u_decod.pc_q_o[7] ),
    .Y(_02005_));
 sky130_fd_sc_hd__and3_1 _06749_ (.A(\u_decod.pc_q_o[6] ),
    .B(\u_decod.pc_q_o[7] ),
    .C(_01917_),
    .X(_02006_));
 sky130_fd_sc_hd__a22o_1 _06750_ (.A1(net39),
    .A2(_01489_),
    .B1(_01490_),
    .B2(net57),
    .X(_02007_));
 sky130_fd_sc_hd__a221o_1 _06751_ (.A1(net62),
    .A2(_01487_),
    .B1(_01488_),
    .B2(net48),
    .C1(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__nand2_1 _06752_ (.A(_01059_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__a22o_1 _06753_ (.A1(_01326_),
    .A2(_01429_),
    .B1(_01435_),
    .B2(_01327_),
    .X(_02010_));
 sky130_fd_sc_hd__a21oi_1 _06754_ (.A1(_01335_),
    .A2(_01432_),
    .B1(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__o311a_1 _06755_ (.A1(_01764_),
    .A2(_02005_),
    .A3(_02006_),
    .B1(_02009_),
    .C1(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__o2111a_1 _06756_ (.A1(_01765_),
    .A2(_01993_),
    .B1(_01998_),
    .C1(_02004_),
    .D1(_02012_),
    .X(_02013_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(_02013_),
    .Y(\u_decod.exe_ff_res_data_i[7] ));
 sky130_fd_sc_hd__a22o_1 _06758_ (.A1(\u_rf.reg11_q[7] ),
    .A2(_01582_),
    .B1(_01634_),
    .B2(\u_rf.reg9_q[7] ),
    .X(_02014_));
 sky130_fd_sc_hd__a221o_1 _06759_ (.A1(\u_rf.reg23_q[7] ),
    .A2(_01612_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[7] ),
    .C1(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a22o_1 _06760_ (.A1(\u_rf.reg16_q[7] ),
    .A2(_01563_),
    .B1(_01651_),
    .B2(\u_rf.reg22_q[7] ),
    .X(_02016_));
 sky130_fd_sc_hd__a221o_1 _06761_ (.A1(\u_rf.reg14_q[7] ),
    .A2(_01657_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[7] ),
    .C1(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__a22o_1 _06762_ (.A1(\u_rf.reg25_q[7] ),
    .A2(_01574_),
    .B1(_01614_),
    .B2(\u_rf.reg31_q[7] ),
    .X(_02018_));
 sky130_fd_sc_hd__a221o_1 _06763_ (.A1(\u_rf.reg12_q[7] ),
    .A2(_01608_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[7] ),
    .C1(_02018_),
    .X(_02019_));
 sky130_fd_sc_hd__a22o_1 _06764_ (.A1(\u_rf.reg5_q[7] ),
    .A2(_01567_),
    .B1(_01620_),
    .B2(\u_rf.reg24_q[7] ),
    .X(_02020_));
 sky130_fd_sc_hd__a221o_1 _06765_ (.A1(\u_rf.reg30_q[7] ),
    .A2(_01579_),
    .B1(_01655_),
    .B2(\u_rf.reg10_q[7] ),
    .C1(_02020_),
    .X(_02021_));
 sky130_fd_sc_hd__or4_1 _06766_ (.A(_02015_),
    .B(_02017_),
    .C(_02019_),
    .D(_02021_),
    .X(_02022_));
 sky130_fd_sc_hd__a22o_1 _06767_ (.A1(\u_rf.reg0_q[7] ),
    .A2(_01516_),
    .B1(_01585_),
    .B2(\u_rf.reg1_q[7] ),
    .X(_02023_));
 sky130_fd_sc_hd__a221o_1 _06768_ (.A1(\u_rf.reg15_q[7] ),
    .A2(_01600_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[7] ),
    .C1(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__a22o_1 _06769_ (.A1(\u_rf.reg26_q[7] ),
    .A2(_01640_),
    .B1(_01643_),
    .B2(\u_rf.reg20_q[7] ),
    .X(_02025_));
 sky130_fd_sc_hd__a221o_1 _06770_ (.A1(\u_rf.reg19_q[7] ),
    .A2(_01594_),
    .B1(_01627_),
    .B2(\u_rf.reg29_q[7] ),
    .C1(_02025_),
    .X(_02026_));
 sky130_fd_sc_hd__a22o_1 _06771_ (.A1(\u_rf.reg18_q[7] ),
    .A2(_01590_),
    .B1(_01623_),
    .B2(\u_rf.reg28_q[7] ),
    .X(_02027_));
 sky130_fd_sc_hd__a221o_1 _06772_ (.A1(\u_rf.reg6_q[7] ),
    .A2(_01554_),
    .B1(_01630_),
    .B2(\u_rf.reg17_q[7] ),
    .C1(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__a22o_1 _06773_ (.A1(\u_rf.reg7_q[7] ),
    .A2(_01559_),
    .B1(_01672_),
    .B2(\u_rf.reg2_q[7] ),
    .X(_02029_));
 sky130_fd_sc_hd__a221o_1 _06774_ (.A1(\u_rf.reg13_q[7] ),
    .A2(_01597_),
    .B1(_01605_),
    .B2(\u_rf.reg3_q[7] ),
    .C1(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__or4_1 _06775_ (.A(_02024_),
    .B(_02026_),
    .C(_02028_),
    .D(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__or2_1 _06776_ (.A(_02022_),
    .B(_02031_),
    .X(_02032_));
 sky130_fd_sc_hd__and2_1 _06777_ (.A(_01679_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__a221o_1 _06778_ (.A1(\u_decod.dec0.funct7[2] ),
    .A2(_01530_),
    .B1(_01549_),
    .B2(\u_decod.rf_ff_res_data_i[7] ),
    .C1(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__a21o_1 _06779_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[7] ),
    .B1(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__nor2_1 _06780_ (.A(_01944_),
    .B(_01990_),
    .Y(_02036_));
 sky130_fd_sc_hd__a21o_1 _06781_ (.A1(_01945_),
    .A2(_02036_),
    .B1(net201),
    .X(_02037_));
 sky130_fd_sc_hd__xnor2_1 _06782_ (.A(_02035_),
    .B(_02037_),
    .Y(\u_decod.rs2_data_nxt[7] ));
 sky130_fd_sc_hd__mux4_1 _06783_ (.A0(\u_decod.rs1_data_q[23] ),
    .A1(_01683_),
    .A2(\u_decod.rs1_data_q[15] ),
    .A3(_01267_),
    .S0(_01445_),
    .S1(_01684_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _06784_ (.A0(_01868_),
    .A1(_02038_),
    .S(_01450_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _06785_ (.A0(_01951_),
    .A1(_02039_),
    .S(_01315_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _06786_ (.A0(_01996_),
    .A1(_02040_),
    .S(_01422_),
    .X(_02041_));
 sky130_fd_sc_hd__o21a_1 _06787_ (.A1(\u_decod.rs1_data_q[8] ),
    .A2(_01445_),
    .B1(_01494_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _06788_ (.A0(_01495_),
    .A1(_02042_),
    .S(_01684_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _06789_ (.A0(_01865_),
    .A1(_02043_),
    .S(_01457_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _06790_ (.A0(_01957_),
    .A1(_02044_),
    .S(_01474_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _06791_ (.A0(_02002_),
    .A1(_02045_),
    .S(_01478_),
    .X(_02046_));
 sky130_fd_sc_hd__a31o_2 _06792_ (.A1(net99),
    .A2(_01064_),
    .A3(_01067_),
    .B1(net100),
    .X(_02047_));
 sky130_fd_sc_hd__and3_1 _06793_ (.A(net99),
    .B(net112),
    .C(_01066_),
    .X(_02048_));
 sky130_fd_sc_hd__buf_2 _06794_ (.A(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__and3b_1 _06795_ (.A_N(\u_decod.unsign_ext_q_o ),
    .B(net62),
    .C(net98),
    .X(_02050_));
 sky130_fd_sc_hd__clkbuf_2 _06796_ (.A(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__a221o_1 _06797_ (.A1(net63),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net49),
    .C1(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__nor2_1 _06798_ (.A(\u_decod.pc_q_o[8] ),
    .B(_02006_),
    .Y(_02053_));
 sky130_fd_sc_hd__and4_2 _06799_ (.A(\u_decod.pc_q_o[6] ),
    .B(\u_decod.pc_q_o[7] ),
    .C(\u_decod.pc_q_o[8] ),
    .D(_01917_),
    .X(_02054_));
 sky130_fd_sc_hd__nand2_1 _06800_ (.A(_01307_),
    .B(_01434_),
    .Y(_02055_));
 sky130_fd_sc_hd__o211a_1 _06801_ (.A1(_01307_),
    .A2(_01763_),
    .B1(_01819_),
    .C1(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__o32a_1 _06802_ (.A1(_01764_),
    .A2(_02053_),
    .A3(_02054_),
    .B1(_02056_),
    .B2(_01339_),
    .X(_02057_));
 sky130_fd_sc_hd__a21bo_1 _06803_ (.A1(_01058_),
    .A2(_02052_),
    .B1_N(_02057_),
    .X(_02058_));
 sky130_fd_sc_hd__o21ai_1 _06804_ (.A1(_01332_),
    .A2(_01336_),
    .B1(_01340_),
    .Y(_02059_));
 sky130_fd_sc_hd__or3_1 _06805_ (.A(_01340_),
    .B(_01332_),
    .C(_01336_),
    .X(_02060_));
 sky130_fd_sc_hd__and3_1 _06806_ (.A(_02059_),
    .B(_01436_),
    .C(_02060_),
    .X(_02061_));
 sky130_fd_sc_hd__a211o_1 _06807_ (.A1(_01504_),
    .A2(_02046_),
    .B1(_02058_),
    .C1(_02061_),
    .X(_02062_));
 sky130_fd_sc_hd__a21oi_1 _06808_ (.A1(_01441_),
    .A2(_02041_),
    .B1(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__inv_2 _06809_ (.A(_02063_),
    .Y(\u_decod.exe_ff_res_data_i[8] ));
 sky130_fd_sc_hd__a22o_1 _06810_ (.A1(\u_rf.reg30_q[8] ),
    .A2(_01578_),
    .B1(_01623_),
    .B2(\u_rf.reg28_q[8] ),
    .X(_02064_));
 sky130_fd_sc_hd__a221o_1 _06811_ (.A1(\u_rf.reg13_q[8] ),
    .A2(_01596_),
    .B1(_01590_),
    .B2(\u_rf.reg18_q[8] ),
    .C1(_02064_),
    .X(_02065_));
 sky130_fd_sc_hd__a22o_1 _06812_ (.A1(\u_rf.reg26_q[8] ),
    .A2(_01640_),
    .B1(_01643_),
    .B2(\u_rf.reg20_q[8] ),
    .X(_02066_));
 sky130_fd_sc_hd__a221o_1 _06813_ (.A1(\u_rf.reg25_q[8] ),
    .A2(_01574_),
    .B1(_01620_),
    .B2(\u_rf.reg24_q[8] ),
    .C1(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__a22o_1 _06814_ (.A1(\u_rf.reg14_q[8] ),
    .A2(_01657_),
    .B1(_01669_),
    .B2(\u_rf.reg27_q[8] ),
    .X(_02068_));
 sky130_fd_sc_hd__a221o_1 _06815_ (.A1(\u_rf.reg29_q[8] ),
    .A2(_01626_),
    .B1(_01637_),
    .B2(\u_rf.reg21_q[8] ),
    .C1(_02068_),
    .X(_02069_));
 sky130_fd_sc_hd__a22o_1 _06816_ (.A1(\u_rf.reg31_q[8] ),
    .A2(_01614_),
    .B1(_01648_),
    .B2(\u_rf.reg4_q[8] ),
    .X(_02070_));
 sky130_fd_sc_hd__a221o_1 _06817_ (.A1(\u_rf.reg12_q[8] ),
    .A2(_01607_),
    .B1(_01672_),
    .B2(\u_rf.reg2_q[8] ),
    .C1(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__or4_1 _06818_ (.A(_02065_),
    .B(_02067_),
    .C(_02069_),
    .D(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__a22o_1 _06819_ (.A1(\u_rf.reg16_q[8] ),
    .A2(_01563_),
    .B1(_01629_),
    .B2(\u_rf.reg17_q[8] ),
    .X(_02073_));
 sky130_fd_sc_hd__a221o_1 _06820_ (.A1(\u_rf.reg5_q[8] ),
    .A2(_01567_),
    .B1(_01593_),
    .B2(\u_rf.reg19_q[8] ),
    .C1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__a22o_1 _06821_ (.A1(\u_rf.reg7_q[8] ),
    .A2(_01559_),
    .B1(_01604_),
    .B2(\u_rf.reg3_q[8] ),
    .X(_02075_));
 sky130_fd_sc_hd__a221o_1 _06822_ (.A1(\u_rf.reg0_q[8] ),
    .A2(_01516_),
    .B1(_01599_),
    .B2(\u_rf.reg15_q[8] ),
    .C1(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__a22o_1 _06823_ (.A1(\u_rf.reg11_q[8] ),
    .A2(_01582_),
    .B1(_01665_),
    .B2(\u_rf.reg8_q[8] ),
    .X(_02077_));
 sky130_fd_sc_hd__a221o_1 _06824_ (.A1(\u_rf.reg1_q[8] ),
    .A2(_01585_),
    .B1(_01634_),
    .B2(\u_rf.reg9_q[8] ),
    .C1(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__a22o_1 _06825_ (.A1(\u_rf.reg6_q[8] ),
    .A2(_01554_),
    .B1(_01651_),
    .B2(\u_rf.reg22_q[8] ),
    .X(_02079_));
 sky130_fd_sc_hd__a221o_1 _06826_ (.A1(\u_rf.reg23_q[8] ),
    .A2(_01611_),
    .B1(_01655_),
    .B2(\u_rf.reg10_q[8] ),
    .C1(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__or4_1 _06827_ (.A(_02074_),
    .B(_02076_),
    .C(_02078_),
    .D(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__o21a_1 _06828_ (.A1(_02072_),
    .A2(_02081_),
    .B1(_01678_),
    .X(_02082_));
 sky130_fd_sc_hd__a221o_1 _06829_ (.A1(\u_decod.dec0.funct7[3] ),
    .A2(_01529_),
    .B1(_01548_),
    .B2(\u_decod.rf_ff_res_data_i[8] ),
    .C1(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a21o_1 _06830_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[8] ),
    .B1(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__a221oi_2 _06831_ (.A1(_01093_),
    .A2(_01090_),
    .B1(_01896_),
    .B2(_01079_),
    .C1(_01237_),
    .Y(_02085_));
 sky130_fd_sc_hd__inv_2 _06832_ (.A(_01895_),
    .Y(_02086_));
 sky130_fd_sc_hd__and2b_1 _06833_ (.A_N(_02035_),
    .B(_02036_),
    .X(_02087_));
 sky130_fd_sc_hd__and4_1 _06834_ (.A(_01804_),
    .B(_02086_),
    .C(_01898_),
    .D(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__buf_2 _06835_ (.A(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__nor2_1 _06836_ (.A(_02085_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__xor2_1 _06837_ (.A(_02084_),
    .B(_02090_),
    .X(\u_decod.rs2_data_nxt[8] ));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_01307_),
    .B(_02059_),
    .Y(_02091_));
 sky130_fd_sc_hd__xnor2_1 _06839_ (.A(_02091_),
    .B(_01337_),
    .Y(_02092_));
 sky130_fd_sc_hd__o211a_1 _06840_ (.A1(\u_decod.rs1_data_q[9] ),
    .A2(_01446_),
    .B1(_01684_),
    .C1(_01753_),
    .X(_02093_));
 sky130_fd_sc_hd__a21o_1 _06841_ (.A1(_01455_),
    .A2(_01704_),
    .B1(_02093_),
    .X(_02094_));
 sky130_fd_sc_hd__mux4_2 _06842_ (.A0(_01824_),
    .A1(_01904_),
    .A2(_02001_),
    .A3(_02094_),
    .S0(_01474_),
    .S1(_01458_),
    .X(_02095_));
 sky130_fd_sc_hd__o21a_1 _06843_ (.A1(\u_decod.rs2_data_q[0] ),
    .A2(_02095_),
    .B1(_01504_),
    .X(_02096_));
 sky130_fd_sc_hd__o21ai_1 _06844_ (.A1(_01478_),
    .A2(_02045_),
    .B1(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__o21a_1 _06845_ (.A1(\u_decod.rs1_data_q[16] ),
    .A2(_01702_),
    .B1(_01703_),
    .X(_02098_));
 sky130_fd_sc_hd__o21a_1 _06846_ (.A1(\u_decod.rs1_data_q[24] ),
    .A2(_01702_),
    .B1(_01703_),
    .X(_02099_));
 sky130_fd_sc_hd__mux2_1 _06847_ (.A0(_02098_),
    .A1(_02099_),
    .S(_01444_),
    .X(_02100_));
 sky130_fd_sc_hd__mux2_1 _06848_ (.A0(_01909_),
    .A1(_02100_),
    .S(_01450_),
    .X(_02101_));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(_01995_),
    .A1(_02101_),
    .S(_01315_),
    .X(_02102_));
 sky130_fd_sc_hd__o21a_1 _06850_ (.A1(_01422_),
    .A2(_02040_),
    .B1(_01441_),
    .X(_02103_));
 sky130_fd_sc_hd__o21ai_1 _06851_ (.A1(_01478_),
    .A2(_02102_),
    .B1(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__a221oi_1 _06852_ (.A1(net64),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net50),
    .C1(_02051_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _06853_ (.A(_01306_),
    .B(_01819_),
    .Y(_02106_));
 sky130_fd_sc_hd__a221oi_2 _06854_ (.A1(_01305_),
    .A2(_01428_),
    .B1(_01434_),
    .B2(_01337_),
    .C1(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__a21oi_1 _06855_ (.A1(\u_decod.pc_q_o[9] ),
    .A2(_02054_),
    .B1(_01764_),
    .Y(_02108_));
 sky130_fd_sc_hd__o21ai_1 _06856_ (.A1(\u_decod.pc_q_o[9] ),
    .A2(_02054_),
    .B1(_02108_),
    .Y(_02109_));
 sky130_fd_sc_hd__o211a_1 _06857_ (.A1(_01057_),
    .A2(_02105_),
    .B1(_02107_),
    .C1(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__o2111a_1 _06858_ (.A1(_01765_),
    .A2(_02092_),
    .B1(_02097_),
    .C1(_02104_),
    .D1(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__inv_2 _06859_ (.A(_02111_),
    .Y(\u_decod.exe_ff_res_data_i[9] ));
 sky130_fd_sc_hd__a22o_1 _06860_ (.A1(\u_rf.reg30_q[9] ),
    .A2(_01578_),
    .B1(_01623_),
    .B2(\u_rf.reg28_q[9] ),
    .X(_02112_));
 sky130_fd_sc_hd__a221o_1 _06861_ (.A1(\u_rf.reg13_q[9] ),
    .A2(_01596_),
    .B1(_01590_),
    .B2(\u_rf.reg18_q[9] ),
    .C1(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__a22o_1 _06862_ (.A1(\u_rf.reg26_q[9] ),
    .A2(_01640_),
    .B1(_01643_),
    .B2(\u_rf.reg20_q[9] ),
    .X(_02114_));
 sky130_fd_sc_hd__a221o_1 _06863_ (.A1(\u_rf.reg25_q[9] ),
    .A2(_01574_),
    .B1(_01620_),
    .B2(\u_rf.reg24_q[9] ),
    .C1(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__a22o_1 _06864_ (.A1(\u_rf.reg14_q[9] ),
    .A2(_01657_),
    .B1(_01669_),
    .B2(\u_rf.reg27_q[9] ),
    .X(_02116_));
 sky130_fd_sc_hd__a221o_1 _06865_ (.A1(\u_rf.reg29_q[9] ),
    .A2(_01626_),
    .B1(_01637_),
    .B2(\u_rf.reg21_q[9] ),
    .C1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__a22o_1 _06866_ (.A1(\u_rf.reg31_q[9] ),
    .A2(_01614_),
    .B1(_01648_),
    .B2(\u_rf.reg4_q[9] ),
    .X(_02118_));
 sky130_fd_sc_hd__a221o_1 _06867_ (.A1(\u_rf.reg12_q[9] ),
    .A2(_01607_),
    .B1(_01672_),
    .B2(\u_rf.reg2_q[9] ),
    .C1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__or4_1 _06868_ (.A(_02113_),
    .B(_02115_),
    .C(_02117_),
    .D(_02119_),
    .X(_02120_));
 sky130_fd_sc_hd__a22o_1 _06869_ (.A1(\u_rf.reg16_q[9] ),
    .A2(_01563_),
    .B1(_01629_),
    .B2(\u_rf.reg17_q[9] ),
    .X(_02121_));
 sky130_fd_sc_hd__a221o_1 _06870_ (.A1(\u_rf.reg5_q[9] ),
    .A2(_01567_),
    .B1(_01593_),
    .B2(\u_rf.reg19_q[9] ),
    .C1(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__a22o_1 _06871_ (.A1(\u_rf.reg7_q[9] ),
    .A2(_01559_),
    .B1(_01604_),
    .B2(\u_rf.reg3_q[9] ),
    .X(_02123_));
 sky130_fd_sc_hd__a221o_1 _06872_ (.A1(\u_rf.reg0_q[9] ),
    .A2(_01516_),
    .B1(_01599_),
    .B2(\u_rf.reg15_q[9] ),
    .C1(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__a22o_1 _06873_ (.A1(\u_rf.reg6_q[9] ),
    .A2(_01554_),
    .B1(_01651_),
    .B2(\u_rf.reg22_q[9] ),
    .X(_02125_));
 sky130_fd_sc_hd__a221o_1 _06874_ (.A1(\u_rf.reg23_q[9] ),
    .A2(_01611_),
    .B1(_01655_),
    .B2(\u_rf.reg10_q[9] ),
    .C1(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__a22o_1 _06875_ (.A1(\u_rf.reg11_q[9] ),
    .A2(_01582_),
    .B1(_01665_),
    .B2(\u_rf.reg8_q[9] ),
    .X(_02127_));
 sky130_fd_sc_hd__a221o_1 _06876_ (.A1(\u_rf.reg1_q[9] ),
    .A2(_01585_),
    .B1(_01634_),
    .B2(\u_rf.reg9_q[9] ),
    .C1(_02127_),
    .X(_02128_));
 sky130_fd_sc_hd__or4_1 _06877_ (.A(_02122_),
    .B(_02124_),
    .C(_02126_),
    .D(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__o21a_1 _06878_ (.A1(_02120_),
    .A2(_02129_),
    .B1(_01678_),
    .X(_02130_));
 sky130_fd_sc_hd__a221o_1 _06879_ (.A1(\u_decod.dec0.funct7[4] ),
    .A2(_01529_),
    .B1(_01548_),
    .B2(\u_decod.rf_ff_res_data_i[9] ),
    .C1(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__a21o_1 _06880_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[9] ),
    .B1(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__o21ai_1 _06881_ (.A1(_02084_),
    .A2(_02090_),
    .B1(_01744_),
    .Y(_02133_));
 sky130_fd_sc_hd__xnor2_1 _06882_ (.A(_02132_),
    .B(_02133_),
    .Y(\u_decod.rs2_data_nxt[9] ));
 sky130_fd_sc_hd__o31ai_2 _06883_ (.A1(_01305_),
    .A2(_01308_),
    .A3(_01341_),
    .B1(_01345_),
    .Y(_02134_));
 sky130_fd_sc_hd__or4_1 _06884_ (.A(_01345_),
    .B(_01305_),
    .C(_01308_),
    .D(_01341_),
    .X(_02135_));
 sky130_fd_sc_hd__buf_2 _06885_ (.A(_01703_),
    .X(_02136_));
 sky130_fd_sc_hd__o21a_1 _06886_ (.A1(\u_decod.rs1_data_q[25] ),
    .A2(_01454_),
    .B1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__mux4_1 _06887_ (.A0(_01949_),
    .A1(_01754_),
    .A2(_01950_),
    .A3(_02137_),
    .S0(_01450_),
    .S1(_01467_),
    .X(_02138_));
 sky130_fd_sc_hd__mux2_1 _06888_ (.A0(_02039_),
    .A1(_02138_),
    .S(_01493_),
    .X(_02139_));
 sky130_fd_sc_hd__mux2_1 _06889_ (.A0(_02102_),
    .A1(_02139_),
    .S(_01422_),
    .X(_02140_));
 sky130_fd_sc_hd__o21a_1 _06890_ (.A1(_01302_),
    .A2(_01702_),
    .B1(_01703_),
    .X(_02141_));
 sky130_fd_sc_hd__mux2_1 _06891_ (.A0(_01748_),
    .A1(_02141_),
    .S(_01685_),
    .X(_02142_));
 sky130_fd_sc_hd__o211a_1 _06892_ (.A1(_01460_),
    .A2(_01955_),
    .B1(_01498_),
    .C1(_01450_),
    .X(_02143_));
 sky130_fd_sc_hd__a21oi_1 _06893_ (.A1(_01458_),
    .A2(_02142_),
    .B1(_02143_),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _06894_ (.A(_01315_),
    .B(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__a211o_1 _06895_ (.A1(_01493_),
    .A2(_02044_),
    .B1(_02145_),
    .C1(\u_decod.rs2_data_q[0] ),
    .X(_02146_));
 sky130_fd_sc_hd__o211a_1 _06896_ (.A1(_01478_),
    .A2(_02095_),
    .B1(_02146_),
    .C1(_01505_),
    .X(_02147_));
 sky130_fd_sc_hd__a221o_1 _06897_ (.A1(net34),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net51),
    .C1(_02051_),
    .X(_02148_));
 sky130_fd_sc_hd__a21oi_1 _06898_ (.A1(\u_decod.pc_q_o[9] ),
    .A2(_02054_),
    .B1(\u_decod.pc_q_o[10] ),
    .Y(_02149_));
 sky130_fd_sc_hd__and3_1 _06899_ (.A(\u_decod.pc_q_o[9] ),
    .B(\u_decod.pc_q_o[10] ),
    .C(_02054_),
    .X(_02150_));
 sky130_fd_sc_hd__nand2_1 _06900_ (.A(_01303_),
    .B(_01434_),
    .Y(_02151_));
 sky130_fd_sc_hd__o211a_1 _06901_ (.A1(_01303_),
    .A2(_01763_),
    .B1(_01819_),
    .C1(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__o32a_1 _06902_ (.A1(_01764_),
    .A2(_02149_),
    .A3(_02150_),
    .B1(_02152_),
    .B2(_01344_),
    .X(_02153_));
 sky130_fd_sc_hd__a21bo_1 _06903_ (.A1(_01058_),
    .A2(_02148_),
    .B1_N(_02153_),
    .X(_02154_));
 sky130_fd_sc_hd__a211o_1 _06904_ (.A1(_01441_),
    .A2(_02140_),
    .B1(_02147_),
    .C1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__a31oi_2 _06905_ (.A1(_02134_),
    .A2(_01437_),
    .A3(_02135_),
    .B1(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__inv_2 _06906_ (.A(_02156_),
    .Y(\u_decod.exe_ff_res_data_i[10] ));
 sky130_fd_sc_hd__a22o_1 _06907_ (.A1(\u_rf.reg6_q[10] ),
    .A2(_01554_),
    .B1(_01651_),
    .B2(\u_rf.reg22_q[10] ),
    .X(_02157_));
 sky130_fd_sc_hd__a221o_1 _06908_ (.A1(\u_rf.reg23_q[10] ),
    .A2(_01611_),
    .B1(_01655_),
    .B2(\u_rf.reg10_q[10] ),
    .C1(_02157_),
    .X(_02158_));
 sky130_fd_sc_hd__a22o_1 _06909_ (.A1(\u_rf.reg11_q[10] ),
    .A2(_01582_),
    .B1(_01665_),
    .B2(\u_rf.reg8_q[10] ),
    .X(_02159_));
 sky130_fd_sc_hd__a221o_1 _06910_ (.A1(\u_rf.reg1_q[10] ),
    .A2(_01585_),
    .B1(_01634_),
    .B2(\u_rf.reg9_q[10] ),
    .C1(_02159_),
    .X(_02160_));
 sky130_fd_sc_hd__a22o_1 _06911_ (.A1(\u_rf.reg7_q[10] ),
    .A2(_01559_),
    .B1(_01604_),
    .B2(\u_rf.reg3_q[10] ),
    .X(_02161_));
 sky130_fd_sc_hd__a221o_1 _06912_ (.A1(\u_rf.reg0_q[10] ),
    .A2(_01516_),
    .B1(_01599_),
    .B2(\u_rf.reg15_q[10] ),
    .C1(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__a22o_1 _06913_ (.A1(\u_rf.reg16_q[10] ),
    .A2(_01563_),
    .B1(_01629_),
    .B2(\u_rf.reg17_q[10] ),
    .X(_02163_));
 sky130_fd_sc_hd__a221o_1 _06914_ (.A1(\u_rf.reg5_q[10] ),
    .A2(_01567_),
    .B1(_01594_),
    .B2(\u_rf.reg19_q[10] ),
    .C1(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__or4_1 _06915_ (.A(_02158_),
    .B(_02160_),
    .C(_02162_),
    .D(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__a22o_1 _06916_ (.A1(\u_rf.reg31_q[10] ),
    .A2(_01614_),
    .B1(_01648_),
    .B2(\u_rf.reg4_q[10] ),
    .X(_02166_));
 sky130_fd_sc_hd__a221o_1 _06917_ (.A1(\u_rf.reg12_q[10] ),
    .A2(_01607_),
    .B1(_01672_),
    .B2(\u_rf.reg2_q[10] ),
    .C1(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__a22o_1 _06918_ (.A1(\u_rf.reg14_q[10] ),
    .A2(_01657_),
    .B1(_01669_),
    .B2(\u_rf.reg27_q[10] ),
    .X(_02168_));
 sky130_fd_sc_hd__a221o_1 _06919_ (.A1(\u_rf.reg29_q[10] ),
    .A2(_01626_),
    .B1(_01637_),
    .B2(\u_rf.reg21_q[10] ),
    .C1(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__a22o_1 _06920_ (.A1(\u_rf.reg30_q[10] ),
    .A2(_01578_),
    .B1(_01623_),
    .B2(\u_rf.reg28_q[10] ),
    .X(_02170_));
 sky130_fd_sc_hd__a221o_1 _06921_ (.A1(\u_rf.reg13_q[10] ),
    .A2(_01596_),
    .B1(_01590_),
    .B2(\u_rf.reg18_q[10] ),
    .C1(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__a22o_1 _06922_ (.A1(\u_rf.reg26_q[10] ),
    .A2(_01640_),
    .B1(_01643_),
    .B2(\u_rf.reg20_q[10] ),
    .X(_02172_));
 sky130_fd_sc_hd__a221o_1 _06923_ (.A1(\u_rf.reg25_q[10] ),
    .A2(_01574_),
    .B1(_01620_),
    .B2(\u_rf.reg24_q[10] ),
    .C1(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__or4_1 _06924_ (.A(_02167_),
    .B(_02169_),
    .C(_02171_),
    .D(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__o21a_1 _06925_ (.A1(_02165_),
    .A2(_02174_),
    .B1(_01678_),
    .X(_02175_));
 sky130_fd_sc_hd__a221o_1 _06926_ (.A1(\u_decod.dec0.funct7[5] ),
    .A2(_01530_),
    .B1(_01548_),
    .B2(\u_decod.rf_ff_res_data_i[10] ),
    .C1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__a21o_1 _06927_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[10] ),
    .B1(_02176_),
    .X(_02177_));
 sky130_fd_sc_hd__or2_1 _06928_ (.A(_02084_),
    .B(_02132_),
    .X(_02178_));
 sky130_fd_sc_hd__a21oi_1 _06929_ (.A1(_01897_),
    .A2(_02178_),
    .B1(_02090_),
    .Y(_02179_));
 sky130_fd_sc_hd__xnor2_1 _06930_ (.A(_02177_),
    .B(_02179_),
    .Y(\u_decod.rs2_data_nxt[10] ));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(_01303_),
    .B(_02134_),
    .Y(_02180_));
 sky130_fd_sc_hd__xor2_1 _06932_ (.A(_02180_),
    .B(_01342_),
    .X(_02181_));
 sky130_fd_sc_hd__a22oi_1 _06933_ (.A1(_01300_),
    .A2(_01429_),
    .B1(_01435_),
    .B2(_01342_),
    .Y(_02182_));
 sky130_fd_sc_hd__a221o_1 _06934_ (.A1(net35),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net52),
    .C1(_02051_),
    .X(_02183_));
 sky130_fd_sc_hd__o21ai_1 _06935_ (.A1(\u_decod.pc_q_o[11] ),
    .A2(_02150_),
    .B1(_01484_),
    .Y(_02184_));
 sky130_fd_sc_hd__and4_2 _06936_ (.A(\u_decod.pc_q_o[9] ),
    .B(\u_decod.pc_q_o[10] ),
    .C(\u_decod.pc_q_o[11] ),
    .D(_02054_),
    .X(_02185_));
 sky130_fd_sc_hd__o2bb2a_1 _06937_ (.A1_N(_01059_),
    .A2_N(_02183_),
    .B1(_02184_),
    .B2(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__o211ai_1 _06938_ (.A1(_01301_),
    .A2(_01820_),
    .B1(_02182_),
    .C1(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__or2_1 _06939_ (.A(_01424_),
    .B(_02139_),
    .X(_02188_));
 sky130_fd_sc_hd__clkbuf_4 _06940_ (.A(_01479_),
    .X(_02189_));
 sky130_fd_sc_hd__o21a_1 _06941_ (.A1(\u_decod.rs1_data_q[18] ),
    .A2(_01454_),
    .B1(_01753_),
    .X(_02190_));
 sky130_fd_sc_hd__o21a_1 _06942_ (.A1(\u_decod.rs1_data_q[26] ),
    .A2(_01454_),
    .B1(_01753_),
    .X(_02191_));
 sky130_fd_sc_hd__mux2_1 _06943_ (.A0(_02190_),
    .A1(_02191_),
    .S(_01455_),
    .X(_02192_));
 sky130_fd_sc_hd__mux2_1 _06944_ (.A0(_01994_),
    .A1(_02192_),
    .S(_01451_),
    .X(_02193_));
 sky130_fd_sc_hd__mux2_1 _06945_ (.A0(_02101_),
    .A1(_02193_),
    .S(_01757_),
    .X(_02194_));
 sky130_fd_sc_hd__or2_1 _06946_ (.A(_02189_),
    .B(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__o211a_1 _06947_ (.A1(\u_decod.rs1_data_q[11] ),
    .A2(_01454_),
    .B1(_01685_),
    .C1(_02136_),
    .X(_02196_));
 sky130_fd_sc_hd__a21o_1 _06948_ (.A1(_01460_),
    .A2(_01823_),
    .B1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__mux4_1 _06949_ (.A0(_01904_),
    .A1(_02001_),
    .A2(_02094_),
    .A3(_02197_),
    .S0(_01475_),
    .S1(_01905_),
    .X(_02198_));
 sky130_fd_sc_hd__a211o_1 _06950_ (.A1(_01757_),
    .A2(_02044_),
    .B1(_02145_),
    .C1(_01479_),
    .X(_02199_));
 sky130_fd_sc_hd__o211a_1 _06951_ (.A1(_01424_),
    .A2(_02198_),
    .B1(_02199_),
    .C1(_01506_),
    .X(_02200_));
 sky130_fd_sc_hd__a31o_1 _06952_ (.A1(_01442_),
    .A2(_02188_),
    .A3(_02195_),
    .B1(_02200_),
    .X(_02201_));
 sky130_fd_sc_hd__a211oi_1 _06953_ (.A1(_01437_),
    .A2(_02181_),
    .B1(_02187_),
    .C1(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__inv_2 _06954_ (.A(_02202_),
    .Y(\u_decod.exe_ff_res_data_i[11] ));
 sky130_fd_sc_hd__o21a_1 _06955_ (.A1(_01227_),
    .A2(_01530_),
    .B1(\u_decod.dec0.funct7[6] ),
    .X(_02203_));
 sky130_fd_sc_hd__a221o_2 _06956_ (.A1(\u_decod.dec0.instr_i[20] ),
    .A2(_01205_),
    .B1(_01241_),
    .B2(\u_decod.dec0.instr_i[7] ),
    .C1(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__a22o_1 _06957_ (.A1(\u_rf.reg13_q[11] ),
    .A2(_01597_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[11] ),
    .X(_02205_));
 sky130_fd_sc_hd__a221o_1 _06958_ (.A1(\u_rf.reg31_q[11] ),
    .A2(_01616_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[11] ),
    .C1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__a22o_1 _06959_ (.A1(\u_rf.reg5_q[11] ),
    .A2(_01568_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[11] ),
    .X(_02207_));
 sky130_fd_sc_hd__a221o_1 _06960_ (.A1(\u_rf.reg28_q[11] ),
    .A2(_01625_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[11] ),
    .C1(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__a22o_1 _06961_ (.A1(\u_rf.reg12_q[11] ),
    .A2(_01608_),
    .B1(_01642_),
    .B2(\u_rf.reg26_q[11] ),
    .X(_02209_));
 sky130_fd_sc_hd__a221o_1 _06962_ (.A1(\u_rf.reg1_q[11] ),
    .A2(_01587_),
    .B1(_01606_),
    .B2(\u_rf.reg3_q[11] ),
    .C1(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__a22o_1 _06963_ (.A1(\u_rf.reg16_q[11] ),
    .A2(_01564_),
    .B1(_01583_),
    .B2(\u_rf.reg11_q[11] ),
    .X(_02211_));
 sky130_fd_sc_hd__a221o_1 _06964_ (.A1(\u_rf.reg7_q[11] ),
    .A2(_01561_),
    .B1(_01595_),
    .B2(\u_rf.reg19_q[11] ),
    .C1(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__or4_1 _06965_ (.A(_02206_),
    .B(_02208_),
    .C(_02210_),
    .D(_02212_),
    .X(_02213_));
 sky130_fd_sc_hd__a22o_1 _06966_ (.A1(\u_rf.reg18_q[11] ),
    .A2(_01591_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[11] ),
    .X(_02214_));
 sky130_fd_sc_hd__a221o_1 _06967_ (.A1(\u_rf.reg25_q[11] ),
    .A2(_01576_),
    .B1(_01580_),
    .B2(\u_rf.reg30_q[11] ),
    .C1(_02214_),
    .X(_02215_));
 sky130_fd_sc_hd__a22o_1 _06968_ (.A1(\u_rf.reg29_q[11] ),
    .A2(_01627_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[11] ),
    .X(_02216_));
 sky130_fd_sc_hd__a221o_1 _06969_ (.A1(\u_rf.reg0_q[11] ),
    .A2(_01663_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[11] ),
    .C1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__a22o_1 _06970_ (.A1(\u_rf.reg17_q[11] ),
    .A2(_01630_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[11] ),
    .X(_02218_));
 sky130_fd_sc_hd__a221o_1 _06971_ (.A1(\u_rf.reg20_q[11] ),
    .A2(_01645_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[11] ),
    .C1(_02218_),
    .X(_02219_));
 sky130_fd_sc_hd__a22o_1 _06972_ (.A1(\u_rf.reg15_q[11] ),
    .A2(_01600_),
    .B1(_01612_),
    .B2(\u_rf.reg23_q[11] ),
    .X(_02220_));
 sky130_fd_sc_hd__a221o_1 _06973_ (.A1(\u_rf.reg6_q[11] ),
    .A2(_01556_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[11] ),
    .C1(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__or4_1 _06974_ (.A(_02215_),
    .B(_02217_),
    .C(_02219_),
    .D(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__o21a_2 _06975_ (.A1(_02213_),
    .A2(_02222_),
    .B1(_01679_),
    .X(_02223_));
 sky130_fd_sc_hd__a221o_1 _06976_ (.A1(\u_decod.rf_ff_res_data_i[11] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02204_),
    .C1(_02223_),
    .X(_02224_));
 sky130_fd_sc_hd__a21o_1 _06977_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[11] ),
    .B1(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__or2_1 _06978_ (.A(_02177_),
    .B(_02178_),
    .X(_02226_));
 sky130_fd_sc_hd__inv_2 _06979_ (.A(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__a31o_1 _06980_ (.A1(_01075_),
    .A2(_01078_),
    .A3(_01084_),
    .B1(_01089_),
    .X(_02228_));
 sky130_fd_sc_hd__a211oi_4 _06981_ (.A1(_01079_),
    .A2(_01250_),
    .B1(_01243_),
    .C1(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__a21o_1 _06982_ (.A1(_02089_),
    .A2(_02227_),
    .B1(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__xnor2_1 _06983_ (.A(_02225_),
    .B(_02230_),
    .Y(\u_decod.rs2_data_nxt[11] ));
 sky130_fd_sc_hd__o31ai_1 _06984_ (.A1(_01300_),
    .A2(_01304_),
    .A3(_01346_),
    .B1(_01350_),
    .Y(_02231_));
 sky130_fd_sc_hd__and2_1 _06985_ (.A(_02231_),
    .B(_01436_),
    .X(_02232_));
 sky130_fd_sc_hd__o41a_1 _06986_ (.A1(_01350_),
    .A2(_01300_),
    .A3(_01304_),
    .A4(_01346_),
    .B1(_02232_),
    .X(_02233_));
 sky130_fd_sc_hd__and2_1 _06987_ (.A(\u_decod.pc_q_o[12] ),
    .B(_02185_),
    .X(_02234_));
 sky130_fd_sc_hd__o21ai_1 _06988_ (.A1(\u_decod.pc_q_o[12] ),
    .A2(_02185_),
    .B1(_01484_),
    .Y(_02235_));
 sky130_fd_sc_hd__o21a_1 _06989_ (.A1(\u_decod.rs1_data_q[19] ),
    .A2(_01454_),
    .B1(_01753_),
    .X(_02236_));
 sky130_fd_sc_hd__o21a_1 _06990_ (.A1(\u_decod.rs1_data_q[27] ),
    .A2(_01454_),
    .B1(_01753_),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _06991_ (.A0(_02236_),
    .A1(_02237_),
    .S(_01455_),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _06992_ (.A0(_02038_),
    .A1(_02238_),
    .S(_01451_),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _06993_ (.A0(_02138_),
    .A1(_02239_),
    .S(_01493_),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _06994_ (.A0(_02194_),
    .A1(_02240_),
    .S(_01423_),
    .X(_02241_));
 sky130_fd_sc_hd__a2bb2o_1 _06995_ (.A1_N(_02234_),
    .A2_N(_02235_),
    .B1(_01442_),
    .B2(_02241_),
    .X(_02242_));
 sky130_fd_sc_hd__a221o_1 _06996_ (.A1(net36),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net53),
    .C1(_02051_),
    .X(_02243_));
 sky130_fd_sc_hd__buf_2 _06997_ (.A(_01697_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _06998_ (.A0(_01763_),
    .A1(_02244_),
    .S(_01298_),
    .X(_02245_));
 sky130_fd_sc_hd__a21oi_1 _06999_ (.A1(_01820_),
    .A2(_02245_),
    .B1(_01349_),
    .Y(_02246_));
 sky130_fd_sc_hd__o21a_1 _07000_ (.A1(\u_decod.rs1_data_q[12] ),
    .A2(_01445_),
    .B1(_01494_),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _07001_ (.A0(_01864_),
    .A1(_02247_),
    .S(_01684_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _07002_ (.A0(_02043_),
    .A1(_02248_),
    .S(_01457_),
    .X(_02249_));
 sky130_fd_sc_hd__inv_2 _07003_ (.A(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__mux2_1 _07004_ (.A0(_02144_),
    .A1(_02250_),
    .S(_01474_),
    .X(_02251_));
 sky130_fd_sc_hd__nand2_1 _07005_ (.A(_01479_),
    .B(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__o211a_1 _07006_ (.A1(_02189_),
    .A2(_02198_),
    .B1(_02252_),
    .C1(_01505_),
    .X(_02253_));
 sky130_fd_sc_hd__a211o_1 _07007_ (.A1(_01059_),
    .A2(_02243_),
    .B1(_02246_),
    .C1(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__or3_1 _07008_ (.A(_02233_),
    .B(_02242_),
    .C(_02254_),
    .X(_02255_));
 sky130_fd_sc_hd__buf_1 _07009_ (.A(_02255_),
    .X(\u_decod.exe_ff_res_data_i[12] ));
 sky130_fd_sc_hd__o21a_4 _07010_ (.A1(_01226_),
    .A2(_01530_),
    .B1(\u_decod.dec0.funct7[6] ),
    .X(_02256_));
 sky130_fd_sc_hd__a21o_1 _07011_ (.A1(\u_decod.dec0.funct3[0] ),
    .A2(_01208_),
    .B1(_02256_),
    .X(_02257_));
 sky130_fd_sc_hd__a22o_1 _07012_ (.A1(\u_rf.reg25_q[12] ),
    .A2(_01575_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[12] ),
    .X(_02258_));
 sky130_fd_sc_hd__a221o_1 _07013_ (.A1(\u_rf.reg15_q[12] ),
    .A2(_01601_),
    .B1(_01609_),
    .B2(\u_rf.reg12_q[12] ),
    .C1(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__a22o_1 _07014_ (.A1(\u_rf.reg7_q[12] ),
    .A2(_01560_),
    .B1(_01642_),
    .B2(\u_rf.reg26_q[12] ),
    .X(_02260_));
 sky130_fd_sc_hd__a221o_1 _07015_ (.A1(\u_rf.reg31_q[12] ),
    .A2(_01616_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[12] ),
    .C1(_02260_),
    .X(_02261_));
 sky130_fd_sc_hd__a22o_1 _07016_ (.A1(\u_rf.reg19_q[12] ),
    .A2(_01594_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[12] ),
    .X(_02262_));
 sky130_fd_sc_hd__a221o_1 _07017_ (.A1(\u_rf.reg0_q[12] ),
    .A2(_01663_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[12] ),
    .C1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__a22o_1 _07018_ (.A1(\u_rf.reg5_q[12] ),
    .A2(_01568_),
    .B1(_01555_),
    .B2(\u_rf.reg6_q[12] ),
    .X(_02264_));
 sky130_fd_sc_hd__a221o_1 _07019_ (.A1(\u_rf.reg3_q[12] ),
    .A2(_01606_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[12] ),
    .C1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__or4_1 _07020_ (.A(_02259_),
    .B(_02261_),
    .C(_02263_),
    .D(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__a22o_1 _07021_ (.A1(\u_rf.reg30_q[12] ),
    .A2(_01579_),
    .B1(_01591_),
    .B2(\u_rf.reg18_q[12] ),
    .X(_02267_));
 sky130_fd_sc_hd__a221o_1 _07022_ (.A1(\u_rf.reg11_q[12] ),
    .A2(_01584_),
    .B1(_01598_),
    .B2(\u_rf.reg13_q[12] ),
    .C1(_02267_),
    .X(_02268_));
 sky130_fd_sc_hd__a22o_1 _07023_ (.A1(\u_rf.reg29_q[12] ),
    .A2(_01627_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[12] ),
    .X(_02269_));
 sky130_fd_sc_hd__a221o_1 _07024_ (.A1(\u_rf.reg17_q[12] ),
    .A2(_01631_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[12] ),
    .C1(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__a22o_1 _07025_ (.A1(\u_rf.reg1_q[12] ),
    .A2(_01586_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[12] ),
    .X(_02271_));
 sky130_fd_sc_hd__a221o_1 _07026_ (.A1(\u_rf.reg16_q[12] ),
    .A2(_01565_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[12] ),
    .C1(_02271_),
    .X(_02272_));
 sky130_fd_sc_hd__a22o_1 _07027_ (.A1(\u_rf.reg23_q[12] ),
    .A2(_01612_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[12] ),
    .X(_02273_));
 sky130_fd_sc_hd__a221o_1 _07028_ (.A1(\u_rf.reg20_q[12] ),
    .A2(_01645_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[12] ),
    .C1(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__or4_1 _07029_ (.A(_02268_),
    .B(_02270_),
    .C(_02272_),
    .D(_02274_),
    .X(_02275_));
 sky130_fd_sc_hd__o21a_2 _07030_ (.A1(_02266_),
    .A2(_02275_),
    .B1(_01679_),
    .X(_02276_));
 sky130_fd_sc_hd__a221o_1 _07031_ (.A1(\u_decod.rf_ff_res_data_i[12] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02257_),
    .C1(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__a21oi_1 _07032_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[12] ),
    .B1(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__or2_1 _07033_ (.A(_02225_),
    .B(_02226_),
    .X(_02279_));
 sky130_fd_sc_hd__a21o_1 _07034_ (.A1(_01897_),
    .A2(_02279_),
    .B1(_02090_),
    .X(_02280_));
 sky130_fd_sc_hd__xnor2_1 _07035_ (.A(_02278_),
    .B(_02280_),
    .Y(\u_decod.rs2_data_nxt[12] ));
 sky130_fd_sc_hd__nand2_1 _07036_ (.A(_01298_),
    .B(_02231_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _07037_ (.A(_02281_),
    .B(_01347_),
    .Y(_02282_));
 sky130_fd_sc_hd__or2_1 _07038_ (.A(_02281_),
    .B(_01347_),
    .X(_02283_));
 sky130_fd_sc_hd__and3_1 _07039_ (.A(\u_decod.pc_q_o[12] ),
    .B(\u_decod.pc_q_o[13] ),
    .C(_02185_),
    .X(_02284_));
 sky130_fd_sc_hd__o21ai_1 _07040_ (.A1(\u_decod.pc_q_o[13] ),
    .A2(_02234_),
    .B1(_01484_),
    .Y(_02285_));
 sky130_fd_sc_hd__o21a_1 _07041_ (.A1(\u_decod.rs1_data_q[20] ),
    .A2(_01454_),
    .B1(_01753_),
    .X(_02286_));
 sky130_fd_sc_hd__o21a_1 _07042_ (.A1(\u_decod.rs1_data_q[28] ),
    .A2(_01446_),
    .B1(_01753_),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _07043_ (.A0(_02286_),
    .A1(_02287_),
    .S(_01455_),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _07044_ (.A0(_02100_),
    .A1(_02288_),
    .S(_01451_),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _07045_ (.A0(_02193_),
    .A1(_02289_),
    .S(_01493_),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(_02240_),
    .A1(_02290_),
    .S(_01422_),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(_02001_),
    .A1(_02197_),
    .S(_01458_),
    .X(_02292_));
 sky130_fd_sc_hd__o211a_1 _07048_ (.A1(\u_decod.rs1_data_q[13] ),
    .A2(_01454_),
    .B1(_01685_),
    .C1(_02136_),
    .X(_02293_));
 sky130_fd_sc_hd__a21o_1 _07049_ (.A1(_01460_),
    .A2(_01903_),
    .B1(_02293_),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _07050_ (.A0(_02094_),
    .A1(_02294_),
    .S(_01458_),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(_02292_),
    .A1(_02295_),
    .S(_01474_),
    .X(_02296_));
 sky130_fd_sc_hd__nand2_1 _07052_ (.A(_01422_),
    .B(_02251_),
    .Y(_02297_));
 sky130_fd_sc_hd__o211a_1 _07053_ (.A1(_01422_),
    .A2(_02296_),
    .B1(_02297_),
    .C1(_01505_),
    .X(_02298_));
 sky130_fd_sc_hd__a221o_1 _07054_ (.A1(net37),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net54),
    .C1(_02051_),
    .X(_02299_));
 sky130_fd_sc_hd__or2_1 _07055_ (.A(_01295_),
    .B(_01697_),
    .X(_02300_));
 sky130_fd_sc_hd__a21oi_1 _07056_ (.A1(_01819_),
    .A2(_02300_),
    .B1(_01296_),
    .Y(_02301_));
 sky130_fd_sc_hd__a221o_1 _07057_ (.A1(_01295_),
    .A2(_01429_),
    .B1(_02299_),
    .B2(_01058_),
    .C1(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__a211o_1 _07058_ (.A1(_01441_),
    .A2(_02291_),
    .B1(_02298_),
    .C1(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__o21bai_1 _07059_ (.A1(_02284_),
    .A2(_02285_),
    .B1_N(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__a31o_1 _07060_ (.A1(_01437_),
    .A2(_02282_),
    .A3(_02283_),
    .B1(_02304_),
    .X(\u_decod.exe_ff_res_data_i[13] ));
 sky130_fd_sc_hd__nor2_1 _07061_ (.A(_01206_),
    .B(_01530_),
    .Y(_02305_));
 sky130_fd_sc_hd__a21oi_2 _07062_ (.A1(\u_decod.dec0.funct3[1] ),
    .A2(_01208_),
    .B1(_02256_),
    .Y(_02306_));
 sky130_fd_sc_hd__clkbuf_8 _07063_ (.A(_01565_),
    .X(_02307_));
 sky130_fd_sc_hd__a22o_1 _07064_ (.A1(\u_rf.reg1_q[13] ),
    .A2(_01587_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[13] ),
    .X(_02308_));
 sky130_fd_sc_hd__a221o_1 _07065_ (.A1(\u_rf.reg16_q[13] ),
    .A2(_02307_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[13] ),
    .C1(_02308_),
    .X(_02309_));
 sky130_fd_sc_hd__a22o_1 _07066_ (.A1(\u_rf.reg25_q[13] ),
    .A2(_01575_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[13] ),
    .X(_02310_));
 sky130_fd_sc_hd__a221o_1 _07067_ (.A1(\u_rf.reg15_q[13] ),
    .A2(_01601_),
    .B1(_01608_),
    .B2(\u_rf.reg12_q[13] ),
    .C1(_02310_),
    .X(_02311_));
 sky130_fd_sc_hd__a22o_1 _07068_ (.A1(\u_rf.reg7_q[13] ),
    .A2(_01560_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[13] ),
    .X(_02312_));
 sky130_fd_sc_hd__a221o_1 _07069_ (.A1(\u_rf.reg31_q[13] ),
    .A2(_01615_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[13] ),
    .C1(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__a22o_1 _07070_ (.A1(\u_rf.reg19_q[13] ),
    .A2(_01594_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[13] ),
    .X(_02314_));
 sky130_fd_sc_hd__a221o_1 _07071_ (.A1(\u_rf.reg0_q[13] ),
    .A2(_01663_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[13] ),
    .C1(_02314_),
    .X(_02315_));
 sky130_fd_sc_hd__a22o_1 _07072_ (.A1(\u_rf.reg5_q[13] ),
    .A2(_01568_),
    .B1(_01555_),
    .B2(\u_rf.reg6_q[13] ),
    .X(_02316_));
 sky130_fd_sc_hd__a221o_1 _07073_ (.A1(\u_rf.reg3_q[13] ),
    .A2(_01606_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[13] ),
    .C1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__or4_1 _07074_ (.A(_02311_),
    .B(_02313_),
    .C(_02315_),
    .D(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__a22o_1 _07075_ (.A1(\u_rf.reg23_q[13] ),
    .A2(_01612_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[13] ),
    .X(_02319_));
 sky130_fd_sc_hd__a221o_1 _07076_ (.A1(\u_rf.reg20_q[13] ),
    .A2(_01645_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[13] ),
    .C1(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__a22o_1 _07077_ (.A1(\u_rf.reg30_q[13] ),
    .A2(_01579_),
    .B1(_01591_),
    .B2(\u_rf.reg18_q[13] ),
    .X(_02321_));
 sky130_fd_sc_hd__a221o_1 _07078_ (.A1(\u_rf.reg11_q[13] ),
    .A2(_01584_),
    .B1(_01598_),
    .B2(\u_rf.reg13_q[13] ),
    .C1(_02321_),
    .X(_02322_));
 sky130_fd_sc_hd__a22o_1 _07079_ (.A1(\u_rf.reg29_q[13] ),
    .A2(_01627_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[13] ),
    .X(_02323_));
 sky130_fd_sc_hd__a221o_1 _07080_ (.A1(\u_rf.reg17_q[13] ),
    .A2(_01631_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[13] ),
    .C1(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__or3_1 _07081_ (.A(_02320_),
    .B(_02322_),
    .C(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__o31a_1 _07082_ (.A1(_02309_),
    .A2(_02318_),
    .A3(_02325_),
    .B1(_01679_),
    .X(_02326_));
 sky130_fd_sc_hd__a221o_1 _07083_ (.A1(\u_decod.rf_ff_res_data_i[13] ),
    .A2(_01549_),
    .B1(\u_decod.exe_ff_res_data_i[13] ),
    .B2(_01713_),
    .C1(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__o21ba_1 _07084_ (.A1(_02305_),
    .A2(_02306_),
    .B1_N(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__o21ba_1 _07085_ (.A1(net199),
    .A2(_02278_),
    .B1_N(_02280_),
    .X(_02329_));
 sky130_fd_sc_hd__xor2_1 _07086_ (.A(_02328_),
    .B(_02329_),
    .X(\u_decod.rs2_data_nxt[13] ));
 sky130_fd_sc_hd__nor4_1 _07087_ (.A(_01355_),
    .B(_01295_),
    .C(_01299_),
    .D(_01351_),
    .Y(_02330_));
 sky130_fd_sc_hd__o31ai_2 _07088_ (.A1(_01295_),
    .A2(_01299_),
    .A3(_01351_),
    .B1(_01355_),
    .Y(_02331_));
 sky130_fd_sc_hd__clkbuf_4 _07089_ (.A(_01437_),
    .X(_02332_));
 sky130_fd_sc_hd__nand2_1 _07090_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__buf_2 _07091_ (.A(_01764_),
    .X(_02334_));
 sky130_fd_sc_hd__and4_1 _07092_ (.A(\u_decod.pc_q_o[12] ),
    .B(\u_decod.pc_q_o[13] ),
    .C(\u_decod.pc_q_o[14] ),
    .D(_02185_),
    .X(_02335_));
 sky130_fd_sc_hd__nor2_1 _07093_ (.A(\u_decod.pc_q_o[14] ),
    .B(_02284_),
    .Y(_02336_));
 sky130_fd_sc_hd__or3_1 _07094_ (.A(_02334_),
    .B(_02335_),
    .C(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__o21a_1 _07095_ (.A1(\u_decod.rs1_data_q[14] ),
    .A2(_01446_),
    .B1(_01753_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _07096_ (.A0(_01955_),
    .A1(_02338_),
    .S(_01685_),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _07097_ (.A0(_02142_),
    .A1(_02339_),
    .S(_01457_),
    .X(_02340_));
 sky130_fd_sc_hd__mux4_2 _07098_ (.A0(_02292_),
    .A1(_02249_),
    .A2(_02295_),
    .A3(_02340_),
    .S0(_01480_),
    .S1(_01477_),
    .X(_02341_));
 sky130_fd_sc_hd__a221o_1 _07099_ (.A1(net38),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net56),
    .C1(_02051_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _07100_ (.A0(_01763_),
    .A1(_02244_),
    .S(_01293_),
    .X(_02343_));
 sky130_fd_sc_hd__a21oi_1 _07101_ (.A1(_01820_),
    .A2(_02343_),
    .B1(_01354_),
    .Y(_02344_));
 sky130_fd_sc_hd__inv_2 _07102_ (.A(_02239_),
    .Y(_02345_));
 sky130_fd_sc_hd__o21a_1 _07103_ (.A1(\u_decod.rs1_data_q[29] ),
    .A2(_01447_),
    .B1(_02136_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _07104_ (.A0(_01950_),
    .A1(_02346_),
    .S(_01467_),
    .X(_02347_));
 sky130_fd_sc_hd__or2_1 _07105_ (.A(_01455_),
    .B(_01754_),
    .X(_02348_));
 sky130_fd_sc_hd__o211a_1 _07106_ (.A1(_01685_),
    .A2(_02137_),
    .B1(_02348_),
    .C1(_01458_),
    .X(_02349_));
 sky130_fd_sc_hd__a21oi_1 _07107_ (.A1(_01464_),
    .A2(_02347_),
    .B1(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__mux2_1 _07108_ (.A0(_02345_),
    .A1(_02350_),
    .S(_01757_),
    .X(_02351_));
 sky130_fd_sc_hd__nand2_1 _07109_ (.A(_01425_),
    .B(_02351_),
    .Y(_02352_));
 sky130_fd_sc_hd__o211a_1 _07110_ (.A1(_01425_),
    .A2(_02290_),
    .B1(_02352_),
    .C1(_01442_),
    .X(_02353_));
 sky130_fd_sc_hd__a211o_1 _07111_ (.A1(net133),
    .A2(_02342_),
    .B1(_02344_),
    .C1(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__a21oi_1 _07112_ (.A1(_01746_),
    .A2(_02341_),
    .B1(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__o211a_1 _07113_ (.A1(_02330_),
    .A2(_02333_),
    .B1(_02337_),
    .C1(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__inv_2 _07114_ (.A(_02356_),
    .Y(\u_decod.exe_ff_res_data_i[14] ));
 sky130_fd_sc_hd__buf_2 _07115_ (.A(_01772_),
    .X(_02357_));
 sky130_fd_sc_hd__clkbuf_4 _07116_ (.A(_01550_),
    .X(_02358_));
 sky130_fd_sc_hd__buf_4 _07117_ (.A(_01680_),
    .X(_02359_));
 sky130_fd_sc_hd__clkbuf_8 _07118_ (.A(_01636_),
    .X(_02360_));
 sky130_fd_sc_hd__a22o_1 _07119_ (.A1(\u_rf.reg19_q[14] ),
    .A2(_01595_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[14] ),
    .X(_02361_));
 sky130_fd_sc_hd__a221o_1 _07120_ (.A1(\u_rf.reg0_q[14] ),
    .A2(_01664_),
    .B1(_02360_),
    .B2(\u_rf.reg9_q[14] ),
    .C1(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__clkbuf_8 _07121_ (.A(_01606_),
    .X(_02363_));
 sky130_fd_sc_hd__clkbuf_8 _07122_ (.A(_01639_),
    .X(_02364_));
 sky130_fd_sc_hd__a22o_1 _07123_ (.A1(\u_rf.reg5_q[14] ),
    .A2(_01569_),
    .B1(_01556_),
    .B2(\u_rf.reg6_q[14] ),
    .X(_02365_));
 sky130_fd_sc_hd__a221o_1 _07124_ (.A1(\u_rf.reg3_q[14] ),
    .A2(_02363_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[14] ),
    .C1(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__clkbuf_8 _07125_ (.A(_01659_),
    .X(_02367_));
 sky130_fd_sc_hd__buf_4 _07126_ (.A(_01642_),
    .X(_02368_));
 sky130_fd_sc_hd__a22o_1 _07127_ (.A1(\u_rf.reg7_q[14] ),
    .A2(_01561_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[14] ),
    .X(_02369_));
 sky130_fd_sc_hd__a221o_1 _07128_ (.A1(\u_rf.reg31_q[14] ),
    .A2(_01777_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[14] ),
    .C1(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__clkbuf_8 _07129_ (.A(_01601_),
    .X(_02371_));
 sky130_fd_sc_hd__a22o_1 _07130_ (.A1(\u_rf.reg25_q[14] ),
    .A2(_01576_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[14] ),
    .X(_02372_));
 sky130_fd_sc_hd__a221o_1 _07131_ (.A1(\u_rf.reg15_q[14] ),
    .A2(_02371_),
    .B1(_01610_),
    .B2(\u_rf.reg12_q[14] ),
    .C1(_02372_),
    .X(_02373_));
 sky130_fd_sc_hd__or4_1 _07132_ (.A(_02362_),
    .B(_02366_),
    .C(_02370_),
    .D(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__buf_4 _07133_ (.A(_01584_),
    .X(_02375_));
 sky130_fd_sc_hd__clkbuf_8 _07134_ (.A(_01598_),
    .X(_02376_));
 sky130_fd_sc_hd__a22o_1 _07135_ (.A1(\u_rf.reg30_q[14] ),
    .A2(_01580_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[14] ),
    .X(_02377_));
 sky130_fd_sc_hd__a221o_1 _07136_ (.A1(\u_rf.reg11_q[14] ),
    .A2(_02375_),
    .B1(_02376_),
    .B2(\u_rf.reg13_q[14] ),
    .C1(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__clkbuf_8 _07137_ (.A(_01631_),
    .X(_02379_));
 sky130_fd_sc_hd__clkbuf_8 _07138_ (.A(_01791_),
    .X(_02380_));
 sky130_fd_sc_hd__a22o_1 _07139_ (.A1(\u_rf.reg29_q[14] ),
    .A2(_01628_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[14] ),
    .X(_02381_));
 sky130_fd_sc_hd__a221o_1 _07140_ (.A1(\u_rf.reg17_q[14] ),
    .A2(_02379_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[14] ),
    .C1(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__a22o_1 _07141_ (.A1(\u_rf.reg1_q[14] ),
    .A2(_01587_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[14] ),
    .X(_02383_));
 sky130_fd_sc_hd__a221o_1 _07142_ (.A1(\u_rf.reg16_q[14] ),
    .A2(_02307_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[14] ),
    .C1(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__clkbuf_8 _07143_ (.A(_01645_),
    .X(_02385_));
 sky130_fd_sc_hd__buf_4 _07144_ (.A(_01671_),
    .X(_02386_));
 sky130_fd_sc_hd__a22o_1 _07145_ (.A1(\u_rf.reg23_q[14] ),
    .A2(_01613_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[14] ),
    .X(_02387_));
 sky130_fd_sc_hd__a221o_1 _07146_ (.A1(\u_rf.reg20_q[14] ),
    .A2(_02385_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[14] ),
    .C1(_02387_),
    .X(_02388_));
 sky130_fd_sc_hd__or4_1 _07147_ (.A(_02378_),
    .B(_02382_),
    .C(_02384_),
    .D(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__or2_1 _07148_ (.A(_02374_),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__a21oi_2 _07149_ (.A1(\u_decod.dec0.funct3[2] ),
    .A2(_01208_),
    .B1(_02256_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _07150_ (.A(_02305_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__a221o_1 _07151_ (.A1(\u_decod.rf_ff_res_data_i[14] ),
    .A2(_02358_),
    .B1(_02359_),
    .B2(_02390_),
    .C1(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__a21o_1 _07152_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[14] ),
    .B1(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__and4b_1 _07153_ (.A_N(_02225_),
    .B(_02227_),
    .C(_02278_),
    .D(_02328_),
    .X(_02395_));
 sky130_fd_sc_hd__a21oi_1 _07154_ (.A1(_02089_),
    .A2(_02395_),
    .B1(net201),
    .Y(_02396_));
 sky130_fd_sc_hd__xor2_1 _07155_ (.A(_02394_),
    .B(_02396_),
    .X(\u_decod.rs2_data_nxt[14] ));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(_01293_),
    .B(_02331_),
    .Y(_02397_));
 sky130_fd_sc_hd__xor2_1 _07157_ (.A(_02397_),
    .B(_01352_),
    .X(_02398_));
 sky130_fd_sc_hd__o211a_1 _07158_ (.A1(_01289_),
    .A2(_01447_),
    .B1(_01685_),
    .C1(_02136_),
    .X(_02399_));
 sky130_fd_sc_hd__a21o_1 _07159_ (.A1(_01467_),
    .A2(_02000_),
    .B1(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _07160_ (.A0(_02197_),
    .A1(_02400_),
    .S(_01905_),
    .X(_02401_));
 sky130_fd_sc_hd__mux4_1 _07161_ (.A0(_02249_),
    .A1(_02295_),
    .A2(_02340_),
    .A3(_02401_),
    .S0(_02189_),
    .S1(_01476_),
    .X(_02402_));
 sky130_fd_sc_hd__o21a_1 _07162_ (.A1(_01371_),
    .A2(_01447_),
    .B1(_02136_),
    .X(_02403_));
 sky130_fd_sc_hd__o21a_1 _07163_ (.A1(\u_decod.rs1_data_q[30] ),
    .A2(_01454_),
    .B1(_02136_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _07164_ (.A0(_02403_),
    .A1(_02404_),
    .S(_01460_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _07165_ (.A0(_02192_),
    .A1(_02405_),
    .S(_01451_),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _07166_ (.A0(_02289_),
    .A1(_02406_),
    .S(_01688_),
    .X(_02407_));
 sky130_fd_sc_hd__o21ai_1 _07167_ (.A1(_01480_),
    .A2(_02407_),
    .B1(_01442_),
    .Y(_02408_));
 sky130_fd_sc_hd__a21oi_1 _07168_ (.A1(_01480_),
    .A2(_02351_),
    .B1(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__a221o_1 _07169_ (.A1(net39),
    .A2(_02047_),
    .B1(_02049_),
    .B2(net57),
    .C1(_02051_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_1 _07170_ (.A(\u_decod.rs2_data_q[15] ),
    .B(_01289_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21oi_1 _07171_ (.A1(_02411_),
    .A2(_01435_),
    .B1(_01432_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _07172_ (.A(_01291_),
    .B(_02412_),
    .Y(_02413_));
 sky130_fd_sc_hd__a221o_1 _07173_ (.A1(_01290_),
    .A2(_01429_),
    .B1(_02410_),
    .B2(_01059_),
    .C1(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__a211o_1 _07174_ (.A1(_01746_),
    .A2(_02402_),
    .B1(_02409_),
    .C1(_02414_),
    .X(_02415_));
 sky130_fd_sc_hd__o21ai_1 _07175_ (.A1(\u_decod.pc_q_o[15] ),
    .A2(_02335_),
    .B1(_01485_),
    .Y(_02416_));
 sky130_fd_sc_hd__a21oi_1 _07176_ (.A1(\u_decod.pc_q_o[15] ),
    .A2(_02335_),
    .B1(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__a211o_1 _07177_ (.A1(_01437_),
    .A2(_02398_),
    .B1(_02415_),
    .C1(_02417_),
    .X(\u_decod.exe_ff_res_data_i[15] ));
 sky130_fd_sc_hd__a21oi_1 _07178_ (.A1(\u_decod.dec0.instr_i[15] ),
    .A2(_01208_),
    .B1(_02256_),
    .Y(_02418_));
 sky130_fd_sc_hd__buf_4 _07179_ (.A(_01625_),
    .X(_02419_));
 sky130_fd_sc_hd__a22o_1 _07180_ (.A1(\u_rf.reg25_q[15] ),
    .A2(_01783_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[15] ),
    .X(_02420_));
 sky130_fd_sc_hd__a221o_1 _07181_ (.A1(\u_rf.reg15_q[15] ),
    .A2(_02371_),
    .B1(_01610_),
    .B2(\u_rf.reg12_q[15] ),
    .C1(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__a22o_1 _07182_ (.A1(\u_rf.reg7_q[15] ),
    .A2(_01561_),
    .B1(_01642_),
    .B2(\u_rf.reg26_q[15] ),
    .X(_02422_));
 sky130_fd_sc_hd__a221o_1 _07183_ (.A1(\u_rf.reg31_q[15] ),
    .A2(_01616_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[15] ),
    .C1(_02422_),
    .X(_02423_));
 sky130_fd_sc_hd__a22o_1 _07184_ (.A1(\u_rf.reg5_q[15] ),
    .A2(_01569_),
    .B1(_01556_),
    .B2(\u_rf.reg6_q[15] ),
    .X(_02424_));
 sky130_fd_sc_hd__a221o_1 _07185_ (.A1(\u_rf.reg3_q[15] ),
    .A2(_02363_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[15] ),
    .C1(_02424_),
    .X(_02425_));
 sky130_fd_sc_hd__a22o_1 _07186_ (.A1(\u_rf.reg19_q[15] ),
    .A2(_01595_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[15] ),
    .X(_02426_));
 sky130_fd_sc_hd__a221o_1 _07187_ (.A1(\u_rf.reg0_q[15] ),
    .A2(_01664_),
    .B1(_02360_),
    .B2(\u_rf.reg9_q[15] ),
    .C1(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__or3_1 _07188_ (.A(_02423_),
    .B(_02425_),
    .C(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__a22o_1 _07189_ (.A1(\u_rf.reg30_q[15] ),
    .A2(_01580_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[15] ),
    .X(_02429_));
 sky130_fd_sc_hd__a221o_1 _07190_ (.A1(\u_rf.reg11_q[15] ),
    .A2(_01584_),
    .B1(_02376_),
    .B2(\u_rf.reg13_q[15] ),
    .C1(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__a22o_1 _07191_ (.A1(\u_rf.reg29_q[15] ),
    .A2(_01628_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[15] ),
    .X(_02431_));
 sky130_fd_sc_hd__a221o_1 _07192_ (.A1(\u_rf.reg17_q[15] ),
    .A2(_02379_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[15] ),
    .C1(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__a22o_1 _07193_ (.A1(\u_rf.reg1_q[15] ),
    .A2(_01587_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[15] ),
    .X(_02433_));
 sky130_fd_sc_hd__a221o_1 _07194_ (.A1(\u_rf.reg16_q[15] ),
    .A2(_02307_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[15] ),
    .C1(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__a22o_1 _07195_ (.A1(\u_rf.reg23_q[15] ),
    .A2(_01613_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[15] ),
    .X(_02435_));
 sky130_fd_sc_hd__a221o_1 _07196_ (.A1(\u_rf.reg20_q[15] ),
    .A2(_02385_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[15] ),
    .C1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__or4_1 _07197_ (.A(_02430_),
    .B(_02432_),
    .C(_02434_),
    .D(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__o31a_2 _07198_ (.A1(_02421_),
    .A2(_02428_),
    .A3(_02437_),
    .B1(_01680_),
    .X(_02438_));
 sky130_fd_sc_hd__a221o_1 _07199_ (.A1(\u_decod.rf_ff_res_data_i[15] ),
    .A2(_01550_),
    .B1(\u_decod.exe_ff_res_data_i[15] ),
    .B2(_01772_),
    .C1(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__o21ba_1 _07200_ (.A1(_02305_),
    .A2(_02418_),
    .B1_N(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__o21a_1 _07201_ (.A1(_02394_),
    .A2(_02396_),
    .B1(_01744_),
    .X(_02441_));
 sky130_fd_sc_hd__xnor2_1 _07202_ (.A(_02440_),
    .B(_02441_),
    .Y(\u_decod.rs2_data_nxt[15] ));
 sky130_fd_sc_hd__or2_1 _07203_ (.A(_01357_),
    .B(_01391_),
    .X(_02442_));
 sky130_fd_sc_hd__o31ai_4 _07204_ (.A1(_01290_),
    .A2(_01294_),
    .A3(_01356_),
    .B1(_01391_),
    .Y(_02443_));
 sky130_fd_sc_hd__and4_1 _07205_ (.A(net99),
    .B(net39),
    .C(_01064_),
    .D(_01067_),
    .X(_02444_));
 sky130_fd_sc_hd__a221o_1 _07206_ (.A1(net98),
    .A2(net62),
    .B1(net57),
    .B2(_02049_),
    .C1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__nand2b_2 _07207_ (.A_N(\u_decod.unsign_ext_q_o ),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(net40),
    .B(net100),
    .Y(_02447_));
 sky130_fd_sc_hd__a21oi_1 _07209_ (.A1(_02446_),
    .A2(_02447_),
    .B1(_01057_),
    .Y(_02448_));
 sky130_fd_sc_hd__mux4_1 _07210_ (.A0(_01388_),
    .A1(\u_decod.rs1_data_q[8] ),
    .A2(_01061_),
    .A3(_01747_),
    .S0(_01455_),
    .S1(_01461_),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _07211_ (.A0(_02248_),
    .A1(_02449_),
    .S(_01458_),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_1 _07212_ (.A0(_02295_),
    .A1(_02340_),
    .A2(_02401_),
    .A3(_02450_),
    .S0(_01478_),
    .S1(_01475_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _07213_ (.A0(_01763_),
    .A1(_02244_),
    .S(_01400_),
    .X(_02452_));
 sky130_fd_sc_hd__a21oi_1 _07214_ (.A1(_01820_),
    .A2(_02452_),
    .B1(_01390_),
    .Y(_02453_));
 sky130_fd_sc_hd__o211a_1 _07215_ (.A1(_01367_),
    .A2(_01447_),
    .B1(_01685_),
    .C1(_02136_),
    .X(_02454_));
 sky130_fd_sc_hd__a31o_1 _07216_ (.A1(_01267_),
    .A2(_01467_),
    .A3(_02136_),
    .B1(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _07217_ (.A0(_02238_),
    .A1(_02455_),
    .S(_01464_),
    .X(_02456_));
 sky130_fd_sc_hd__nor2_1 _07218_ (.A(_01688_),
    .B(_02350_),
    .Y(_02457_));
 sky130_fd_sc_hd__a211o_1 _07219_ (.A1(_01688_),
    .A2(_02456_),
    .B1(_02457_),
    .C1(_01478_),
    .X(_02458_));
 sky130_fd_sc_hd__o211a_1 _07220_ (.A1(_01422_),
    .A2(_02407_),
    .B1(_02458_),
    .C1(_01441_),
    .X(_02459_));
 sky130_fd_sc_hd__a211o_1 _07221_ (.A1(_01505_),
    .A2(_02451_),
    .B1(_02453_),
    .C1(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__and3_1 _07222_ (.A(\u_decod.pc_q_o[15] ),
    .B(\u_decod.pc_q_o[16] ),
    .C(_02335_),
    .X(_02461_));
 sky130_fd_sc_hd__a21oi_1 _07223_ (.A1(\u_decod.pc_q_o[15] ),
    .A2(_02335_),
    .B1(\u_decod.pc_q_o[16] ),
    .Y(_02462_));
 sky130_fd_sc_hd__or3_1 _07224_ (.A(_01764_),
    .B(_02461_),
    .C(_02462_),
    .X(_02463_));
 sky130_fd_sc_hd__or3b_1 _07225_ (.A(_02448_),
    .B(_02460_),
    .C_N(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__a31o_1 _07226_ (.A1(_01437_),
    .A2(_02442_),
    .A3(_02443_),
    .B1(_02464_),
    .X(\u_decod.exe_ff_res_data_i[16] ));
 sky130_fd_sc_hd__a21o_1 _07227_ (.A1(\u_decod.dec0.instr_i[16] ),
    .A2(_01208_),
    .B1(_02256_),
    .X(_02465_));
 sky130_fd_sc_hd__a22o_1 _07228_ (.A1(\u_rf.reg1_q[16] ),
    .A2(_01587_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[16] ),
    .X(_02466_));
 sky130_fd_sc_hd__a221o_1 _07229_ (.A1(\u_rf.reg16_q[16] ),
    .A2(_01565_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[16] ),
    .C1(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__a22o_1 _07230_ (.A1(\u_rf.reg25_q[16] ),
    .A2(_01575_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[16] ),
    .X(_02468_));
 sky130_fd_sc_hd__a221o_1 _07231_ (.A1(\u_rf.reg15_q[16] ),
    .A2(_01600_),
    .B1(_01608_),
    .B2(\u_rf.reg12_q[16] ),
    .C1(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__a22o_1 _07232_ (.A1(\u_rf.reg7_q[16] ),
    .A2(_01560_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[16] ),
    .X(_02470_));
 sky130_fd_sc_hd__a221o_1 _07233_ (.A1(\u_rf.reg31_q[16] ),
    .A2(_01615_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[16] ),
    .C1(_02470_),
    .X(_02471_));
 sky130_fd_sc_hd__a22o_1 _07234_ (.A1(\u_rf.reg19_q[16] ),
    .A2(_01594_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[16] ),
    .X(_02472_));
 sky130_fd_sc_hd__a221o_1 _07235_ (.A1(\u_rf.reg0_q[16] ),
    .A2(_01662_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[16] ),
    .C1(_02472_),
    .X(_02473_));
 sky130_fd_sc_hd__a22o_1 _07236_ (.A1(\u_rf.reg5_q[16] ),
    .A2(_01568_),
    .B1(_01555_),
    .B2(\u_rf.reg6_q[16] ),
    .X(_02474_));
 sky130_fd_sc_hd__a221o_1 _07237_ (.A1(\u_rf.reg3_q[16] ),
    .A2(_01605_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[16] ),
    .C1(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__or4_1 _07238_ (.A(_02469_),
    .B(_02471_),
    .C(_02473_),
    .D(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__a22o_1 _07239_ (.A1(\u_rf.reg23_q[16] ),
    .A2(_01612_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[16] ),
    .X(_02477_));
 sky130_fd_sc_hd__a221o_1 _07240_ (.A1(\u_rf.reg20_q[16] ),
    .A2(_01644_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[16] ),
    .C1(_02477_),
    .X(_02478_));
 sky130_fd_sc_hd__a22o_1 _07241_ (.A1(\u_rf.reg30_q[16] ),
    .A2(_01579_),
    .B1(_01591_),
    .B2(\u_rf.reg18_q[16] ),
    .X(_02479_));
 sky130_fd_sc_hd__a221o_1 _07242_ (.A1(\u_rf.reg11_q[16] ),
    .A2(_01583_),
    .B1(_01597_),
    .B2(\u_rf.reg13_q[16] ),
    .C1(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__a22o_1 _07243_ (.A1(\u_rf.reg29_q[16] ),
    .A2(_01627_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[16] ),
    .X(_02481_));
 sky130_fd_sc_hd__a221o_1 _07244_ (.A1(\u_rf.reg17_q[16] ),
    .A2(_01630_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[16] ),
    .C1(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__or3_1 _07245_ (.A(_02478_),
    .B(_02480_),
    .C(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__o31a_2 _07246_ (.A1(_02467_),
    .A2(_02476_),
    .A3(_02483_),
    .B1(_01679_),
    .X(_02484_));
 sky130_fd_sc_hd__a221o_1 _07247_ (.A1(\u_decod.rf_ff_res_data_i[16] ),
    .A2(_01549_),
    .B1(_01714_),
    .B2(_02465_),
    .C1(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__a21o_1 _07248_ (.A1(_01713_),
    .A2(\u_decod.exe_ff_res_data_i[16] ),
    .B1(_02485_),
    .X(_02486_));
 sky130_fd_sc_hd__and3b_1 _07249_ (.A_N(_02394_),
    .B(_02395_),
    .C(_02440_),
    .X(_02487_));
 sky130_fd_sc_hd__nand2_1 _07250_ (.A(_02089_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nand2_1 _07251_ (.A(_01897_),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__xnor2_1 _07252_ (.A(_02486_),
    .B(_02489_),
    .Y(\u_decod.rs2_data_nxt[16] ));
 sky130_fd_sc_hd__a21o_1 _07253_ (.A1(_01400_),
    .A2(_02443_),
    .B1(_01383_),
    .X(_02490_));
 sky130_fd_sc_hd__nand3_1 _07254_ (.A(_01400_),
    .B(_01383_),
    .C(_02443_),
    .Y(_02491_));
 sky130_fd_sc_hd__a21bo_1 _07255_ (.A1(net100),
    .A2(net41),
    .B1_N(_02446_),
    .X(_02492_));
 sky130_fd_sc_hd__o21a_1 _07256_ (.A1(_01468_),
    .A2(_02099_),
    .B1(_01498_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _07257_ (.A0(_02288_),
    .A1(_02493_),
    .S(_01472_),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(_02406_),
    .A1(_02494_),
    .S(_01757_),
    .X(_02495_));
 sky130_fd_sc_hd__a211o_1 _07259_ (.A1(_01757_),
    .A2(_02456_),
    .B1(_02457_),
    .C1(_01423_),
    .X(_02496_));
 sky130_fd_sc_hd__o211a_1 _07260_ (.A1(_02189_),
    .A2(_02495_),
    .B1(_02496_),
    .C1(_01441_),
    .X(_02497_));
 sky130_fd_sc_hd__mux4_2 _07261_ (.A0(_01380_),
    .A1(\u_decod.rs1_data_q[9] ),
    .A2(\u_decod.rs1_data_q[1] ),
    .A3(_01747_),
    .S0(_01460_),
    .S1(_01461_),
    .X(_02498_));
 sky130_fd_sc_hd__mux4_2 _07262_ (.A0(_02197_),
    .A1(_02294_),
    .A2(_02400_),
    .A3(_02498_),
    .S0(_01474_),
    .S1(_01905_),
    .X(_02499_));
 sky130_fd_sc_hd__and2_1 _07263_ (.A(_01493_),
    .B(_02340_),
    .X(_02500_));
 sky130_fd_sc_hd__a211o_1 _07264_ (.A1(_01475_),
    .A2(_02450_),
    .B1(_02500_),
    .C1(_01478_),
    .X(_02501_));
 sky130_fd_sc_hd__o211a_1 _07265_ (.A1(_01422_),
    .A2(_02499_),
    .B1(_02501_),
    .C1(_01505_),
    .X(_02502_));
 sky130_fd_sc_hd__a2bb2o_1 _07266_ (.A1_N(_01383_),
    .A2_N(_02244_),
    .B1(_01431_),
    .B2(_01382_),
    .X(_02503_));
 sky130_fd_sc_hd__a311o_1 _07267_ (.A1(\u_decod.rs2_data_q[17] ),
    .A2(_01380_),
    .A3(_01429_),
    .B1(_02502_),
    .C1(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__a211o_1 _07268_ (.A1(_01059_),
    .A2(_02492_),
    .B1(_02497_),
    .C1(_02504_),
    .X(_02505_));
 sky130_fd_sc_hd__and4_1 _07269_ (.A(\u_decod.pc_q_o[15] ),
    .B(\u_decod.pc_q_o[16] ),
    .C(\u_decod.pc_q_o[17] ),
    .D(_02335_),
    .X(_02506_));
 sky130_fd_sc_hd__nor2_1 _07270_ (.A(_02334_),
    .B(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__o21a_1 _07271_ (.A1(\u_decod.pc_q_o[17] ),
    .A2(_02461_),
    .B1(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__a311o_1 _07272_ (.A1(_01437_),
    .A2(_02490_),
    .A3(_02491_),
    .B1(_02505_),
    .C1(_02508_),
    .X(\u_decod.exe_ff_res_data_i[17] ));
 sky130_fd_sc_hd__a21o_1 _07273_ (.A1(\u_decod.dec0.instr_i[17] ),
    .A2(_01208_),
    .B1(_02256_),
    .X(_02509_));
 sky130_fd_sc_hd__a22o_1 _07274_ (.A1(\u_rf.reg1_q[17] ),
    .A2(_01587_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[17] ),
    .X(_02510_));
 sky130_fd_sc_hd__a221o_1 _07275_ (.A1(\u_rf.reg16_q[17] ),
    .A2(_01565_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[17] ),
    .C1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__a22o_1 _07276_ (.A1(\u_rf.reg25_q[17] ),
    .A2(_01575_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[17] ),
    .X(_02512_));
 sky130_fd_sc_hd__a221o_1 _07277_ (.A1(\u_rf.reg15_q[17] ),
    .A2(_01600_),
    .B1(_01608_),
    .B2(\u_rf.reg12_q[17] ),
    .C1(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__a22o_1 _07278_ (.A1(\u_rf.reg7_q[17] ),
    .A2(_01560_),
    .B1(_01641_),
    .B2(\u_rf.reg26_q[17] ),
    .X(_02514_));
 sky130_fd_sc_hd__a221o_1 _07279_ (.A1(\u_rf.reg31_q[17] ),
    .A2(_01615_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[17] ),
    .C1(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__a22o_1 _07280_ (.A1(\u_rf.reg19_q[17] ),
    .A2(_01594_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[17] ),
    .X(_02516_));
 sky130_fd_sc_hd__a221o_1 _07281_ (.A1(\u_rf.reg0_q[17] ),
    .A2(_01662_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[17] ),
    .C1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__a22o_1 _07282_ (.A1(\u_rf.reg5_q[17] ),
    .A2(_01568_),
    .B1(_01555_),
    .B2(\u_rf.reg6_q[17] ),
    .X(_02518_));
 sky130_fd_sc_hd__a221o_1 _07283_ (.A1(\u_rf.reg3_q[17] ),
    .A2(_01605_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[17] ),
    .C1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__or4_1 _07284_ (.A(_02513_),
    .B(_02515_),
    .C(_02517_),
    .D(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a22o_1 _07285_ (.A1(\u_rf.reg23_q[17] ),
    .A2(_01612_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[17] ),
    .X(_02521_));
 sky130_fd_sc_hd__a221o_1 _07286_ (.A1(\u_rf.reg20_q[17] ),
    .A2(_01644_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[17] ),
    .C1(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__a22o_1 _07287_ (.A1(\u_rf.reg30_q[17] ),
    .A2(_01579_),
    .B1(_01591_),
    .B2(\u_rf.reg18_q[17] ),
    .X(_02523_));
 sky130_fd_sc_hd__a221o_1 _07288_ (.A1(\u_rf.reg11_q[17] ),
    .A2(_01583_),
    .B1(_01598_),
    .B2(\u_rf.reg13_q[17] ),
    .C1(_02523_),
    .X(_02524_));
 sky130_fd_sc_hd__a22o_1 _07289_ (.A1(\u_rf.reg29_q[17] ),
    .A2(_01627_),
    .B1(_01652_),
    .B2(\u_rf.reg22_q[17] ),
    .X(_02525_));
 sky130_fd_sc_hd__a221o_1 _07290_ (.A1(\u_rf.reg17_q[17] ),
    .A2(_01630_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[17] ),
    .C1(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__or3_1 _07291_ (.A(_02522_),
    .B(_02524_),
    .C(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__o31a_1 _07292_ (.A1(_02511_),
    .A2(_02520_),
    .A3(_02527_),
    .B1(_01679_),
    .X(_02528_));
 sky130_fd_sc_hd__a221o_1 _07293_ (.A1(\u_decod.rf_ff_res_data_i[17] ),
    .A2(_01549_),
    .B1(_01773_),
    .B2(_02509_),
    .C1(_02528_),
    .X(_02529_));
 sky130_fd_sc_hd__a21o_1 _07294_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[17] ),
    .B1(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__o21ai_1 _07295_ (.A1(_02486_),
    .A2(_02488_),
    .B1(_01744_),
    .Y(_02531_));
 sky130_fd_sc_hd__xnor2_1 _07296_ (.A(_02530_),
    .B(_02531_),
    .Y(\u_decod.rs2_data_nxt[17] ));
 sky130_fd_sc_hd__a31o_1 _07297_ (.A1(_01381_),
    .A2(_01400_),
    .A3(_02443_),
    .B1(_01401_),
    .X(_02532_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(_01387_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__a311o_1 _07299_ (.A1(_01381_),
    .A2(_01400_),
    .A3(_02443_),
    .B1(_01387_),
    .C1(_01401_),
    .X(_02534_));
 sky130_fd_sc_hd__mux4_1 _07300_ (.A0(_01950_),
    .A1(_02137_),
    .A2(_02346_),
    .A3(_01747_),
    .S0(_01464_),
    .S1(_01468_),
    .X(_02535_));
 sky130_fd_sc_hd__mux2_1 _07301_ (.A0(_02456_),
    .A1(_02535_),
    .S(_01757_),
    .X(_02536_));
 sky130_fd_sc_hd__mux2_1 _07302_ (.A0(_02495_),
    .A1(_02536_),
    .S(_01425_),
    .X(_02537_));
 sky130_fd_sc_hd__nand2_1 _07303_ (.A(net100),
    .B(net42),
    .Y(_02538_));
 sky130_fd_sc_hd__a21oi_1 _07304_ (.A1(_02446_),
    .A2(_02538_),
    .B1(_01057_),
    .Y(_02539_));
 sky130_fd_sc_hd__mux4_1 _07305_ (.A0(_01384_),
    .A1(_01302_),
    .A2(\u_decod.rs1_data_q[2] ),
    .A3(_01747_),
    .S0(_01455_),
    .S1(_01447_),
    .X(_02540_));
 sky130_fd_sc_hd__mux2_1 _07306_ (.A0(_02339_),
    .A1(_02540_),
    .S(_01458_),
    .X(_02541_));
 sky130_fd_sc_hd__or2_1 _07307_ (.A(_01688_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__o21ai_1 _07308_ (.A1(_01475_),
    .A2(_02450_),
    .B1(_02542_),
    .Y(_02543_));
 sky130_fd_sc_hd__nand2_1 _07309_ (.A(_02189_),
    .B(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__o211a_1 _07310_ (.A1(_02189_),
    .A2(_02499_),
    .B1(_02544_),
    .C1(_01505_),
    .X(_02545_));
 sky130_fd_sc_hd__a2bb2o_1 _07311_ (.A1_N(_01387_),
    .A2_N(_02244_),
    .B1(_01432_),
    .B2(_01385_),
    .X(_02546_));
 sky130_fd_sc_hd__a2111o_1 _07312_ (.A1(_01403_),
    .A2(_01429_),
    .B1(_02539_),
    .C1(_02545_),
    .D1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__a21oi_1 _07313_ (.A1(\u_decod.pc_q_o[18] ),
    .A2(_02506_),
    .B1(_02334_),
    .Y(_02548_));
 sky130_fd_sc_hd__o21a_1 _07314_ (.A1(\u_decod.pc_q_o[18] ),
    .A2(_02506_),
    .B1(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__a211o_1 _07315_ (.A1(_01443_),
    .A2(_02537_),
    .B1(_02547_),
    .C1(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__a31o_1 _07316_ (.A1(_02332_),
    .A2(_02533_),
    .A3(_02534_),
    .B1(_02550_),
    .X(\u_decod.exe_ff_res_data_i[18] ));
 sky130_fd_sc_hd__a21o_1 _07317_ (.A1(\u_decod.dec0.instr_i[18] ),
    .A2(_01208_),
    .B1(_02256_),
    .X(_02551_));
 sky130_fd_sc_hd__a22o_1 _07318_ (.A1(\u_rf.reg5_q[18] ),
    .A2(_01568_),
    .B1(_01556_),
    .B2(\u_rf.reg6_q[18] ),
    .X(_02552_));
 sky130_fd_sc_hd__a221o_1 _07319_ (.A1(\u_rf.reg3_q[18] ),
    .A2(_01606_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[18] ),
    .C1(_02552_),
    .X(_02553_));
 sky130_fd_sc_hd__a22o_1 _07320_ (.A1(\u_rf.reg0_q[18] ),
    .A2(_01662_),
    .B1(_01635_),
    .B2(\u_rf.reg9_q[18] ),
    .X(_02554_));
 sky130_fd_sc_hd__a221o_1 _07321_ (.A1(\u_rf.reg19_q[18] ),
    .A2(_01595_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[18] ),
    .C1(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__a22o_1 _07322_ (.A1(\u_rf.reg25_q[18] ),
    .A2(_01576_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[18] ),
    .X(_02556_));
 sky130_fd_sc_hd__a221o_1 _07323_ (.A1(\u_rf.reg15_q[18] ),
    .A2(_01601_),
    .B1(_01609_),
    .B2(\u_rf.reg12_q[18] ),
    .C1(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__a22o_1 _07324_ (.A1(\u_rf.reg7_q[18] ),
    .A2(_01561_),
    .B1(_01642_),
    .B2(\u_rf.reg26_q[18] ),
    .X(_02558_));
 sky130_fd_sc_hd__a221o_1 _07325_ (.A1(\u_rf.reg31_q[18] ),
    .A2(_01616_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[18] ),
    .C1(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__or4_1 _07326_ (.A(_02553_),
    .B(_02555_),
    .C(_02557_),
    .D(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__a22o_1 _07327_ (.A1(\u_rf.reg29_q[18] ),
    .A2(_01627_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[18] ),
    .X(_02561_));
 sky130_fd_sc_hd__a221o_1 _07328_ (.A1(\u_rf.reg17_q[18] ),
    .A2(_01631_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[18] ),
    .C1(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__a22o_1 _07329_ (.A1(\u_rf.reg30_q[18] ),
    .A2(_01580_),
    .B1(_01591_),
    .B2(\u_rf.reg18_q[18] ),
    .X(_02563_));
 sky130_fd_sc_hd__a221o_1 _07330_ (.A1(\u_rf.reg11_q[18] ),
    .A2(_01584_),
    .B1(_01598_),
    .B2(\u_rf.reg13_q[18] ),
    .C1(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__a22o_1 _07331_ (.A1(\u_rf.reg23_q[18] ),
    .A2(_01613_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[18] ),
    .X(_02565_));
 sky130_fd_sc_hd__a221o_1 _07332_ (.A1(\u_rf.reg20_q[18] ),
    .A2(_01645_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[18] ),
    .C1(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__a22o_1 _07333_ (.A1(\u_rf.reg1_q[18] ),
    .A2(_01586_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[18] ),
    .X(_02567_));
 sky130_fd_sc_hd__a221o_1 _07334_ (.A1(\u_rf.reg16_q[18] ),
    .A2(_01565_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[18] ),
    .C1(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__or4_1 _07335_ (.A(_02562_),
    .B(_02564_),
    .C(_02566_),
    .D(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__o21a_2 _07336_ (.A1(_02560_),
    .A2(_02569_),
    .B1(_01680_),
    .X(_02570_));
 sky130_fd_sc_hd__a221o_1 _07337_ (.A1(\u_decod.rf_ff_res_data_i[18] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02551_),
    .C1(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__a21oi_1 _07338_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[18] ),
    .B1(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_1 _07339_ (.A(_02486_),
    .B(_02530_),
    .Y(_02573_));
 sky130_fd_sc_hd__o21ai_1 _07340_ (.A1(net199),
    .A2(_02573_),
    .B1(_02489_),
    .Y(_02574_));
 sky130_fd_sc_hd__xnor2_1 _07341_ (.A(_02572_),
    .B(_02574_),
    .Y(\u_decod.rs2_data_nxt[18] ));
 sky130_fd_sc_hd__a21oi_1 _07342_ (.A1(_01386_),
    .A2(_02534_),
    .B1(_01379_),
    .Y(_02575_));
 sky130_fd_sc_hd__a31o_1 _07343_ (.A1(_01386_),
    .A2(_01379_),
    .A3(_02534_),
    .B1(_01765_),
    .X(_02576_));
 sky130_fd_sc_hd__a21oi_1 _07344_ (.A1(\u_decod.pc_q_o[18] ),
    .A2(_02506_),
    .B1(\u_decod.pc_q_o[19] ),
    .Y(_02577_));
 sky130_fd_sc_hd__and3_1 _07345_ (.A(\u_decod.pc_q_o[18] ),
    .B(\u_decod.pc_q_o[19] ),
    .C(_02506_),
    .X(_02578_));
 sky130_fd_sc_hd__o21a_1 _07346_ (.A1(_01468_),
    .A2(_02191_),
    .B1(_01498_),
    .X(_02579_));
 sky130_fd_sc_hd__mux2_1 _07347_ (.A0(_02405_),
    .A1(_02579_),
    .S(_01472_),
    .X(_02580_));
 sky130_fd_sc_hd__mux2_1 _07348_ (.A0(_02494_),
    .A1(_02580_),
    .S(_01757_),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _07349_ (.A0(_02536_),
    .A1(_02581_),
    .S(_01424_),
    .X(_02582_));
 sky130_fd_sc_hd__a21bo_1 _07350_ (.A1(net100),
    .A2(net43),
    .B1_N(_02446_),
    .X(_02583_));
 sky130_fd_sc_hd__mux4_1 _07351_ (.A0(_01376_),
    .A1(\u_decod.rs1_data_q[11] ),
    .A2(\u_decod.rs1_data_q[3] ),
    .A3(_01747_),
    .S0(_01467_),
    .S1(_01461_),
    .X(_02584_));
 sky130_fd_sc_hd__mux4_1 _07352_ (.A0(_02294_),
    .A1(_02400_),
    .A2(_02498_),
    .A3(_02584_),
    .S0(_01475_),
    .S1(_01905_),
    .X(_02585_));
 sky130_fd_sc_hd__nand2_1 _07353_ (.A(_01423_),
    .B(_02543_),
    .Y(_02586_));
 sky130_fd_sc_hd__o211a_1 _07354_ (.A1(_01423_),
    .A2(_02585_),
    .B1(_02586_),
    .C1(_01505_),
    .X(_02587_));
 sky130_fd_sc_hd__and2_1 _07355_ (.A(_01377_),
    .B(_01378_),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _07356_ (.A1(_01377_),
    .A2(_01431_),
    .B1(_01434_),
    .B2(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__a31o_1 _07357_ (.A1(\u_decod.rs2_data_q[19] ),
    .A2(_01376_),
    .A3(_01429_),
    .B1(_02589_),
    .X(_02590_));
 sky130_fd_sc_hd__a211o_1 _07358_ (.A1(_01059_),
    .A2(_02583_),
    .B1(_02587_),
    .C1(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__a21oi_2 _07359_ (.A1(_01443_),
    .A2(_02582_),
    .B1(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__o31a_1 _07360_ (.A1(_02334_),
    .A2(_02577_),
    .A3(_02578_),
    .B1(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__o21ai_2 _07361_ (.A1(_02575_),
    .A2(_02576_),
    .B1(_02593_),
    .Y(\u_decod.exe_ff_res_data_i[19] ));
 sky130_fd_sc_hd__a21o_1 _07362_ (.A1(\u_decod.dec0.instr_i[19] ),
    .A2(_01208_),
    .B1(_02256_),
    .X(_02594_));
 sky130_fd_sc_hd__a22o_1 _07363_ (.A1(\u_rf.reg2_q[19] ),
    .A2(_01673_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[19] ),
    .X(_02595_));
 sky130_fd_sc_hd__a221o_1 _07364_ (.A1(\u_rf.reg30_q[19] ),
    .A2(_01580_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[19] ),
    .C1(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__a22o_1 _07365_ (.A1(\u_rf.reg31_q[19] ),
    .A2(_01615_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[19] ),
    .X(_02597_));
 sky130_fd_sc_hd__a221o_1 _07366_ (.A1(\u_rf.reg28_q[19] ),
    .A2(_01625_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[19] ),
    .C1(_02597_),
    .X(_02598_));
 sky130_fd_sc_hd__a22o_1 _07367_ (.A1(\u_rf.reg16_q[19] ),
    .A2(_01564_),
    .B1(_01670_),
    .B2(\u_rf.reg27_q[19] ),
    .X(_02599_));
 sky130_fd_sc_hd__a221o_1 _07368_ (.A1(\u_rf.reg23_q[19] ),
    .A2(_01613_),
    .B1(_01609_),
    .B2(\u_rf.reg12_q[19] ),
    .C1(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__a22o_1 _07369_ (.A1(\u_rf.reg11_q[19] ),
    .A2(_01583_),
    .B1(_01642_),
    .B2(\u_rf.reg26_q[19] ),
    .X(_02601_));
 sky130_fd_sc_hd__a221o_1 _07370_ (.A1(\u_rf.reg5_q[19] ),
    .A2(_01569_),
    .B1(_01562_),
    .B2(\u_rf.reg7_q[19] ),
    .C1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__or4_1 _07371_ (.A(_02596_),
    .B(_02598_),
    .C(_02600_),
    .D(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__clkbuf_8 _07372_ (.A(_01586_),
    .X(_02604_));
 sky130_fd_sc_hd__a22o_1 _07373_ (.A1(\u_rf.reg0_q[19] ),
    .A2(_01662_),
    .B1(_01597_),
    .B2(\u_rf.reg13_q[19] ),
    .X(_02605_));
 sky130_fd_sc_hd__a221o_1 _07374_ (.A1(\u_rf.reg1_q[19] ),
    .A2(_02604_),
    .B1(_01576_),
    .B2(\u_rf.reg25_q[19] ),
    .C1(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__a22o_1 _07375_ (.A1(\u_rf.reg15_q[19] ),
    .A2(_01600_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[19] ),
    .X(_02607_));
 sky130_fd_sc_hd__a221o_1 _07376_ (.A1(\u_rf.reg29_q[19] ),
    .A2(_01628_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[19] ),
    .C1(_02607_),
    .X(_02608_));
 sky130_fd_sc_hd__a22o_1 _07377_ (.A1(\u_rf.reg6_q[19] ),
    .A2(_01556_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[19] ),
    .X(_02609_));
 sky130_fd_sc_hd__a221o_1 _07378_ (.A1(\u_rf.reg18_q[19] ),
    .A2(_01592_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[19] ),
    .C1(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__a22o_1 _07379_ (.A1(\u_rf.reg3_q[19] ),
    .A2(_01605_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[19] ),
    .X(_02611_));
 sky130_fd_sc_hd__a221o_1 _07380_ (.A1(\u_rf.reg19_q[19] ),
    .A2(_01595_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[19] ),
    .C1(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__or4_1 _07381_ (.A(_02606_),
    .B(_02608_),
    .C(_02610_),
    .D(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__o21a_2 _07382_ (.A1(_02603_),
    .A2(_02613_),
    .B1(_01680_),
    .X(_02614_));
 sky130_fd_sc_hd__a221o_1 _07383_ (.A1(\u_decod.rf_ff_res_data_i[19] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02594_),
    .C1(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__a21oi_1 _07384_ (.A1(_01772_),
    .A2(\u_decod.exe_ff_res_data_i[19] ),
    .B1(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__a31o_1 _07385_ (.A1(_02489_),
    .A2(_02572_),
    .A3(_02573_),
    .B1(net199),
    .X(_02617_));
 sky130_fd_sc_hd__xor2_1 _07386_ (.A(_02616_),
    .B(_02617_),
    .X(\u_decod.rs2_data_nxt[19] ));
 sky130_fd_sc_hd__clkbuf_2 _07387_ (.A(_02446_),
    .X(_02618_));
 sky130_fd_sc_hd__buf_2 _07388_ (.A(net100),
    .X(_02619_));
 sky130_fd_sc_hd__nand2_1 _07389_ (.A(_02619_),
    .B(net45),
    .Y(_02620_));
 sky130_fd_sc_hd__clkbuf_4 _07390_ (.A(_01057_),
    .X(_02621_));
 sky130_fd_sc_hd__a21oi_1 _07391_ (.A1(_02618_),
    .A2(_02620_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21a_1 _07392_ (.A1(_01468_),
    .A2(_02237_),
    .B1(_01498_),
    .X(_02623_));
 sky130_fd_sc_hd__mux2_1 _07393_ (.A0(_02455_),
    .A1(_02623_),
    .S(_01472_),
    .X(_02624_));
 sky130_fd_sc_hd__mux2_1 _07394_ (.A0(_02535_),
    .A1(_02624_),
    .S(_01757_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(_02581_),
    .A1(_02625_),
    .S(_01424_),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _07396_ (.A0(_01763_),
    .A1(_02244_),
    .S(_01395_),
    .X(_02627_));
 sky130_fd_sc_hd__a21oi_1 _07397_ (.A1(_01820_),
    .A2(_02627_),
    .B1(_01365_),
    .Y(_02628_));
 sky130_fd_sc_hd__mux4_1 _07398_ (.A0(_01363_),
    .A1(_01297_),
    .A2(\u_decod.rs1_data_q[4] ),
    .A3(_01747_),
    .S0(_01460_),
    .S1(_01461_),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _07399_ (.A0(_02449_),
    .A1(_02629_),
    .S(_01905_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _07400_ (.A0(_02541_),
    .A1(_02630_),
    .S(_01475_),
    .X(_02631_));
 sky130_fd_sc_hd__or2_1 _07401_ (.A(_01423_),
    .B(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__o211a_1 _07402_ (.A1(_02189_),
    .A2(_02585_),
    .B1(_02632_),
    .C1(_01506_),
    .X(_02633_));
 sky130_fd_sc_hd__a211o_1 _07403_ (.A1(_01442_),
    .A2(_02626_),
    .B1(_02628_),
    .C1(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__a311o_1 _07404_ (.A1(_02411_),
    .A2(_01293_),
    .A3(_02331_),
    .B1(_01392_),
    .C1(_01291_),
    .X(_02635_));
 sky130_fd_sc_hd__and3_1 _07405_ (.A(_01366_),
    .B(_01405_),
    .C(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__a21oi_1 _07406_ (.A1(_01405_),
    .A2(_02635_),
    .B1(_01366_),
    .Y(_02637_));
 sky130_fd_sc_hd__and2_1 _07407_ (.A(\u_decod.pc_q_o[20] ),
    .B(_02578_),
    .X(_02638_));
 sky130_fd_sc_hd__nor2_1 _07408_ (.A(\u_decod.pc_q_o[20] ),
    .B(_02578_),
    .Y(_02639_));
 sky130_fd_sc_hd__or3_1 _07409_ (.A(_01764_),
    .B(_02638_),
    .C(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__o31a_1 _07410_ (.A1(_01765_),
    .A2(_02636_),
    .A3(_02637_),
    .B1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__or3b_1 _07411_ (.A(_02622_),
    .B(_02634_),
    .C_N(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _07412_ (.A(_02642_),
    .X(\u_decod.exe_ff_res_data_i[20] ));
 sky130_fd_sc_hd__or2_1 _07413_ (.A(_01226_),
    .B(_01715_),
    .X(_02643_));
 sky130_fd_sc_hd__clkbuf_2 _07414_ (.A(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__and2_1 _07415_ (.A(\u_decod.dec0.funct7[6] ),
    .B(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__buf_2 _07416_ (.A(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__a21o_1 _07417_ (.A1(\u_decod.dec0.instr_i[20] ),
    .A2(_01206_),
    .B1(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__a22o_1 _07418_ (.A1(\u_rf.reg27_q[20] ),
    .A2(_01671_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[20] ),
    .X(_02648_));
 sky130_fd_sc_hd__a221o_1 _07419_ (.A1(\u_rf.reg13_q[20] ),
    .A2(_01598_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[20] ),
    .C1(_02648_),
    .X(_02649_));
 sky130_fd_sc_hd__a22o_1 _07420_ (.A1(\u_rf.reg31_q[20] ),
    .A2(_01616_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[20] ),
    .X(_02650_));
 sky130_fd_sc_hd__a221o_1 _07421_ (.A1(\u_rf.reg12_q[20] ),
    .A2(_01609_),
    .B1(_01650_),
    .B2(\u_rf.reg4_q[20] ),
    .C1(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__buf_4 _07422_ (.A(_01613_),
    .X(_02652_));
 sky130_fd_sc_hd__a22o_1 _07423_ (.A1(\u_rf.reg6_q[20] ),
    .A2(_01556_),
    .B1(_01584_),
    .B2(\u_rf.reg11_q[20] ),
    .X(_02653_));
 sky130_fd_sc_hd__a221o_1 _07424_ (.A1(\u_rf.reg23_q[20] ),
    .A2(_02652_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[20] ),
    .C1(_02653_),
    .X(_02654_));
 sky130_fd_sc_hd__a22o_1 _07425_ (.A1(\u_rf.reg30_q[20] ),
    .A2(_01580_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[20] ),
    .X(_02655_));
 sky130_fd_sc_hd__a221o_1 _07426_ (.A1(\u_rf.reg9_q[20] ),
    .A2(_01636_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[20] ),
    .C1(_02655_),
    .X(_02656_));
 sky130_fd_sc_hd__or4_1 _07427_ (.A(_02649_),
    .B(_02651_),
    .C(_02654_),
    .D(_02656_),
    .X(_02657_));
 sky130_fd_sc_hd__a22o_1 _07428_ (.A1(\u_rf.reg26_q[20] ),
    .A2(_01642_),
    .B1(_01645_),
    .B2(\u_rf.reg20_q[20] ),
    .X(_02658_));
 sky130_fd_sc_hd__a221o_1 _07429_ (.A1(\u_rf.reg25_q[20] ),
    .A2(_01576_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[20] ),
    .C1(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__a22o_1 _07430_ (.A1(\u_rf.reg1_q[20] ),
    .A2(_01587_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[20] ),
    .X(_02660_));
 sky130_fd_sc_hd__a221o_1 _07431_ (.A1(\u_rf.reg29_q[20] ),
    .A2(_01628_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[20] ),
    .C1(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__a22o_1 _07432_ (.A1(\u_rf.reg7_q[20] ),
    .A2(_01561_),
    .B1(_01606_),
    .B2(\u_rf.reg3_q[20] ),
    .X(_02662_));
 sky130_fd_sc_hd__a221o_1 _07433_ (.A1(\u_rf.reg0_q[20] ),
    .A2(_01663_),
    .B1(_02371_),
    .B2(\u_rf.reg15_q[20] ),
    .C1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__buf_4 _07434_ (.A(_01569_),
    .X(_02664_));
 sky130_fd_sc_hd__clkbuf_8 _07435_ (.A(_01595_),
    .X(_02665_));
 sky130_fd_sc_hd__a22o_1 _07436_ (.A1(\u_rf.reg16_q[20] ),
    .A2(_01565_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[20] ),
    .X(_02666_));
 sky130_fd_sc_hd__a221o_1 _07437_ (.A1(\u_rf.reg5_q[20] ),
    .A2(_02664_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[20] ),
    .C1(_02666_),
    .X(_02667_));
 sky130_fd_sc_hd__or4_1 _07438_ (.A(_02659_),
    .B(_02661_),
    .C(_02663_),
    .D(_02667_),
    .X(_02668_));
 sky130_fd_sc_hd__o21a_1 _07439_ (.A1(_02657_),
    .A2(_02668_),
    .B1(_01680_),
    .X(_02669_));
 sky130_fd_sc_hd__a221o_1 _07440_ (.A1(\u_decod.rf_ff_res_data_i[20] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02647_),
    .C1(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__a21o_1 _07441_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[20] ),
    .B1(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__and3_1 _07442_ (.A(_02572_),
    .B(_02573_),
    .C(_02616_),
    .X(_02672_));
 sky130_fd_sc_hd__a31o_1 _07443_ (.A1(_02089_),
    .A2(_02487_),
    .A3(_02672_),
    .B1(net199),
    .X(_02673_));
 sky130_fd_sc_hd__xnor2_1 _07444_ (.A(_02671_),
    .B(_02673_),
    .Y(\u_decod.rs2_data_nxt[20] ));
 sky130_fd_sc_hd__a21o_1 _07445_ (.A1(_01405_),
    .A2(_02635_),
    .B1(_01366_),
    .X(_02674_));
 sky130_fd_sc_hd__a21o_1 _07446_ (.A1(_01395_),
    .A2(_02674_),
    .B1(_01362_),
    .X(_02675_));
 sky130_fd_sc_hd__o31a_1 _07447_ (.A1(_01364_),
    .A2(_01361_),
    .A3(_02637_),
    .B1(_02332_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(\u_decod.pc_q_o[21] ),
    .B(_02638_),
    .Y(_02677_));
 sky130_fd_sc_hd__or2_1 _07449_ (.A(\u_decod.pc_q_o[21] ),
    .B(_02638_),
    .X(_02678_));
 sky130_fd_sc_hd__o21a_1 _07450_ (.A1(_01468_),
    .A2(_02287_),
    .B1(_01498_),
    .X(_02679_));
 sky130_fd_sc_hd__mux2_1 _07451_ (.A0(_02493_),
    .A1(_02679_),
    .S(_01472_),
    .X(_02680_));
 sky130_fd_sc_hd__buf_2 _07452_ (.A(_01757_),
    .X(_02681_));
 sky130_fd_sc_hd__mux2_1 _07453_ (.A0(_02580_),
    .A1(_02680_),
    .S(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__mux2_1 _07454_ (.A0(_02625_),
    .A1(_02682_),
    .S(_01425_),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_1 _07455_ (.A0(_01358_),
    .A1(\u_decod.rs1_data_q[13] ),
    .A2(\u_decod.rs1_data_q[5] ),
    .A3(_01747_),
    .S0(_01468_),
    .S1(_01461_),
    .X(_02684_));
 sky130_fd_sc_hd__buf_2 _07456_ (.A(_01905_),
    .X(_02685_));
 sky130_fd_sc_hd__mux4_1 _07457_ (.A0(_02400_),
    .A1(_02498_),
    .A2(_02584_),
    .A3(_02684_),
    .S0(_01475_),
    .S1(_02685_),
    .X(_02686_));
 sky130_fd_sc_hd__mux2_1 _07458_ (.A0(_02631_),
    .A1(_02686_),
    .S(_02189_),
    .X(_02687_));
 sky130_fd_sc_hd__and3_1 _07459_ (.A(\u_decod.rs2_data_q[21] ),
    .B(_01358_),
    .C(\u_decod.instr_operation_q[1] ),
    .X(_02688_));
 sky130_fd_sc_hd__a221o_1 _07460_ (.A1(_01430_),
    .A2(_01360_),
    .B1(_01361_),
    .B2(\u_decod.instr_operation_q[3] ),
    .C1(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__a22o_1 _07461_ (.A1(_01506_),
    .A2(_02687_),
    .B1(_02689_),
    .B2(_01260_),
    .X(_02690_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(_02619_),
    .B(net46),
    .Y(_02691_));
 sky130_fd_sc_hd__a21oi_1 _07463_ (.A1(_02618_),
    .A2(_02691_),
    .B1(_02621_),
    .Y(_02692_));
 sky130_fd_sc_hd__a211o_1 _07464_ (.A1(_01443_),
    .A2(_02683_),
    .B1(_02690_),
    .C1(_02692_),
    .X(_02693_));
 sky130_fd_sc_hd__a31o_1 _07465_ (.A1(_01485_),
    .A2(_02677_),
    .A3(_02678_),
    .B1(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__a21oi_2 _07466_ (.A1(_02675_),
    .A2(_02676_),
    .B1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__inv_2 _07467_ (.A(_02695_),
    .Y(\u_decod.exe_ff_res_data_i[21] ));
 sky130_fd_sc_hd__a21o_1 _07468_ (.A1(\u_decod.dec0.instr_i[21] ),
    .A2(_01206_),
    .B1(_02645_),
    .X(_02696_));
 sky130_fd_sc_hd__buf_4 _07469_ (.A(_01650_),
    .X(_02697_));
 sky130_fd_sc_hd__a22o_1 _07470_ (.A1(\u_rf.reg30_q[21] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[21] ),
    .X(_02698_));
 sky130_fd_sc_hd__a221o_1 _07471_ (.A1(\u_rf.reg31_q[21] ),
    .A2(_01777_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[21] ),
    .C1(_02698_),
    .X(_02699_));
 sky130_fd_sc_hd__a22o_1 _07472_ (.A1(\u_rf.reg12_q[21] ),
    .A2(_01609_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[21] ),
    .X(_02700_));
 sky130_fd_sc_hd__a221o_1 _07473_ (.A1(\u_rf.reg9_q[21] ),
    .A2(_01636_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[21] ),
    .C1(_02700_),
    .X(_02701_));
 sky130_fd_sc_hd__a22o_1 _07474_ (.A1(\u_rf.reg6_q[21] ),
    .A2(_01556_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[21] ),
    .X(_02702_));
 sky130_fd_sc_hd__a221o_1 _07475_ (.A1(\u_rf.reg11_q[21] ),
    .A2(_01584_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[21] ),
    .C1(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__a22o_1 _07476_ (.A1(\u_rf.reg23_q[21] ),
    .A2(_01613_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[21] ),
    .X(_02704_));
 sky130_fd_sc_hd__a221o_1 _07477_ (.A1(\u_rf.reg13_q[21] ),
    .A2(_01598_),
    .B1(_01592_),
    .B2(\u_rf.reg18_q[21] ),
    .C1(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__or3_1 _07478_ (.A(_02701_),
    .B(_02703_),
    .C(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__a22o_1 _07479_ (.A1(\u_rf.reg16_q[21] ),
    .A2(_01564_),
    .B1(_01630_),
    .B2(\u_rf.reg17_q[21] ),
    .X(_02707_));
 sky130_fd_sc_hd__a221o_1 _07480_ (.A1(\u_rf.reg5_q[21] ),
    .A2(_01569_),
    .B1(_01595_),
    .B2(\u_rf.reg19_q[21] ),
    .C1(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__a22o_1 _07481_ (.A1(\u_rf.reg7_q[21] ),
    .A2(_01561_),
    .B1(_01605_),
    .B2(\u_rf.reg3_q[21] ),
    .X(_02709_));
 sky130_fd_sc_hd__a221o_1 _07482_ (.A1(\u_rf.reg0_q[21] ),
    .A2(_01663_),
    .B1(_01601_),
    .B2(\u_rf.reg15_q[21] ),
    .C1(_02709_),
    .X(_02710_));
 sky130_fd_sc_hd__a22o_1 _07483_ (.A1(\u_rf.reg26_q[21] ),
    .A2(_01642_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[21] ),
    .X(_02711_));
 sky130_fd_sc_hd__a221o_1 _07484_ (.A1(\u_rf.reg25_q[21] ),
    .A2(_01576_),
    .B1(_01622_),
    .B2(\u_rf.reg24_q[21] ),
    .C1(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(\u_rf.reg1_q[21] ),
    .A2(_01587_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[21] ),
    .X(_02713_));
 sky130_fd_sc_hd__a221o_1 _07486_ (.A1(\u_rf.reg29_q[21] ),
    .A2(_01628_),
    .B1(_01639_),
    .B2(\u_rf.reg21_q[21] ),
    .C1(_02713_),
    .X(_02714_));
 sky130_fd_sc_hd__or4_1 _07487_ (.A(_02708_),
    .B(_02710_),
    .C(_02712_),
    .D(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__o31a_1 _07488_ (.A1(_02699_),
    .A2(_02706_),
    .A3(_02715_),
    .B1(_01680_),
    .X(_02716_));
 sky130_fd_sc_hd__a221o_1 _07489_ (.A1(\u_decod.rf_ff_res_data_i[21] ),
    .A2(_01550_),
    .B1(_01773_),
    .B2(_02696_),
    .C1(_02716_),
    .X(_02717_));
 sky130_fd_sc_hd__o21bai_2 _07490_ (.A1(_01528_),
    .A2(_02695_),
    .B1_N(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__a21bo_1 _07491_ (.A1(_01897_),
    .A2(_02671_),
    .B1_N(_02673_),
    .X(_02719_));
 sky130_fd_sc_hd__xor2_1 _07492_ (.A(_02718_),
    .B(_02719_),
    .X(\u_decod.rs2_data_nxt[21] ));
 sky130_fd_sc_hd__inv_2 _07493_ (.A(\u_decod.pc_q_o[22] ),
    .Y(_02720_));
 sky130_fd_sc_hd__a31o_1 _07494_ (.A1(\u_decod.pc_q_o[21] ),
    .A2(\u_decod.pc_q_o[22] ),
    .A3(_02638_),
    .B1(_02334_),
    .X(_02721_));
 sky130_fd_sc_hd__a21oi_1 _07495_ (.A1(_02720_),
    .A2(_02677_),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__buf_2 _07496_ (.A(_01425_),
    .X(_02723_));
 sky130_fd_sc_hd__inv_2 _07497_ (.A(_02624_),
    .Y(_02724_));
 sky130_fd_sc_hd__o21a_1 _07498_ (.A1(_01469_),
    .A2(_02346_),
    .B1(_01498_),
    .X(_02725_));
 sky130_fd_sc_hd__o211a_1 _07499_ (.A1(_01469_),
    .A2(_02137_),
    .B1(_01498_),
    .C1(_01905_),
    .X(_02726_));
 sky130_fd_sc_hd__a21oi_1 _07500_ (.A1(_01472_),
    .A2(_02725_),
    .B1(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__mux2_1 _07501_ (.A0(_02724_),
    .A1(_02727_),
    .S(_02681_),
    .X(_02728_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(_01425_),
    .B(_02728_),
    .Y(_02729_));
 sky130_fd_sc_hd__o211a_1 _07503_ (.A1(_02723_),
    .A2(_02682_),
    .B1(_02729_),
    .C1(_01443_),
    .X(_02730_));
 sky130_fd_sc_hd__a21bo_1 _07504_ (.A1(_02619_),
    .A2(net47),
    .B1_N(_02446_),
    .X(_02731_));
 sky130_fd_sc_hd__mux4_1 _07505_ (.A0(_01371_),
    .A1(_01292_),
    .A2(\u_decod.rs1_data_q[6] ),
    .A3(_01747_),
    .S0(_01467_),
    .S1(_01461_),
    .X(_02732_));
 sky130_fd_sc_hd__mux2_1 _07506_ (.A0(_02540_),
    .A1(_02732_),
    .S(_01905_),
    .X(_02733_));
 sky130_fd_sc_hd__mux2_1 _07507_ (.A0(_02630_),
    .A1(_02733_),
    .S(_01476_),
    .X(_02734_));
 sky130_fd_sc_hd__mux2_1 _07508_ (.A0(_02686_),
    .A1(_02734_),
    .S(_01480_),
    .X(_02735_));
 sky130_fd_sc_hd__a22o_1 _07509_ (.A1(net133),
    .A2(_02731_),
    .B1(_02735_),
    .B2(_01746_),
    .X(_02736_));
 sky130_fd_sc_hd__a221o_1 _07510_ (.A1(_01372_),
    .A2(_01373_),
    .B1(_01361_),
    .B2(_02637_),
    .C1(_01397_),
    .X(_02737_));
 sky130_fd_sc_hd__a311o_1 _07511_ (.A1(_01359_),
    .A2(_01395_),
    .A3(_02674_),
    .B1(_01374_),
    .C1(_01396_),
    .X(_02738_));
 sky130_fd_sc_hd__nor2_1 _07512_ (.A(_01374_),
    .B(_02244_),
    .Y(_02739_));
 sky130_fd_sc_hd__a221o_1 _07513_ (.A1(_01398_),
    .A2(_01429_),
    .B1(_01432_),
    .B2(_01372_),
    .C1(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__a31o_1 _07514_ (.A1(_01437_),
    .A2(_02737_),
    .A3(_02738_),
    .B1(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__or4_1 _07515_ (.A(_02722_),
    .B(_02730_),
    .C(_02736_),
    .D(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__buf_1 _07516_ (.A(_02742_),
    .X(\u_decod.exe_ff_res_data_i[22] ));
 sky130_fd_sc_hd__clkbuf_4 _07517_ (.A(_01773_),
    .X(_02743_));
 sky130_fd_sc_hd__a21o_1 _07518_ (.A1(\u_decod.dec0.instr_i[22] ),
    .A2(_01206_),
    .B1(_02646_),
    .X(_02744_));
 sky130_fd_sc_hd__a22o_1 _07519_ (.A1(\u_rf.reg0_q[22] ),
    .A2(_01663_),
    .B1(_01616_),
    .B2(\u_rf.reg31_q[22] ),
    .X(_02745_));
 sky130_fd_sc_hd__a221o_1 _07520_ (.A1(\u_rf.reg3_q[22] ),
    .A2(_02363_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[22] ),
    .C1(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a22o_1 _07521_ (.A1(\u_rf.reg25_q[22] ),
    .A2(_01576_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[22] ),
    .X(_02747_));
 sky130_fd_sc_hd__a221o_1 _07522_ (.A1(\u_rf.reg6_q[22] ),
    .A2(_01557_),
    .B1(_02604_),
    .B2(\u_rf.reg1_q[22] ),
    .C1(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__a22o_1 _07523_ (.A1(\u_rf.reg15_q[22] ),
    .A2(_01601_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[22] ),
    .X(_02749_));
 sky130_fd_sc_hd__a221o_1 _07524_ (.A1(\u_rf.reg14_q[22] ),
    .A2(_02367_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[22] ),
    .C1(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__a22o_1 _07525_ (.A1(\u_rf.reg7_q[22] ),
    .A2(_01562_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[22] ),
    .X(_02751_));
 sky130_fd_sc_hd__a221o_1 _07526_ (.A1(\u_rf.reg16_q[22] ),
    .A2(_02307_),
    .B1(_02376_),
    .B2(\u_rf.reg13_q[22] ),
    .C1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__or4_1 _07527_ (.A(_02746_),
    .B(_02748_),
    .C(_02750_),
    .D(_02752_),
    .X(_02753_));
 sky130_fd_sc_hd__a22o_1 _07528_ (.A1(\u_rf.reg12_q[22] ),
    .A2(_01609_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[22] ),
    .X(_02754_));
 sky130_fd_sc_hd__a221o_1 _07529_ (.A1(\u_rf.reg9_q[22] ),
    .A2(_02360_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[22] ),
    .C1(_02754_),
    .X(_02755_));
 sky130_fd_sc_hd__a22o_1 _07530_ (.A1(\u_rf.reg27_q[22] ),
    .A2(_01671_),
    .B1(_01667_),
    .B2(\u_rf.reg8_q[22] ),
    .X(_02756_));
 sky130_fd_sc_hd__a221o_1 _07531_ (.A1(\u_rf.reg5_q[22] ),
    .A2(_02664_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[22] ),
    .C1(_02756_),
    .X(_02757_));
 sky130_fd_sc_hd__a22o_1 _07532_ (.A1(\u_rf.reg30_q[22] ),
    .A2(_01580_),
    .B1(_01625_),
    .B2(\u_rf.reg28_q[22] ),
    .X(_02758_));
 sky130_fd_sc_hd__a221o_1 _07533_ (.A1(\u_rf.reg17_q[22] ),
    .A2(_02379_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[22] ),
    .C1(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__a22o_1 _07534_ (.A1(\u_rf.reg24_q[22] ),
    .A2(_01622_),
    .B1(_01780_),
    .B2(\u_rf.reg29_q[22] ),
    .X(_02760_));
 sky130_fd_sc_hd__a221o_1 _07535_ (.A1(\u_rf.reg18_q[22] ),
    .A2(_01787_),
    .B1(_02652_),
    .B2(\u_rf.reg23_q[22] ),
    .C1(_02760_),
    .X(_02761_));
 sky130_fd_sc_hd__or4_1 _07536_ (.A(_02755_),
    .B(_02757_),
    .C(_02759_),
    .D(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__o21a_1 _07537_ (.A1(_02753_),
    .A2(_02762_),
    .B1(_02359_),
    .X(_02763_));
 sky130_fd_sc_hd__a221o_1 _07538_ (.A1(\u_decod.rf_ff_res_data_i[22] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_02744_),
    .C1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__a21oi_1 _07539_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[22] ),
    .B1(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _07540_ (.A(_02671_),
    .B(_02718_),
    .Y(_02766_));
 sky130_fd_sc_hd__a41o_1 _07541_ (.A1(_02089_),
    .A2(_02487_),
    .A3(_02672_),
    .A4(_02766_),
    .B1(net200),
    .X(_02767_));
 sky130_fd_sc_hd__and2_1 _07542_ (.A(_02765_),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__nor2_1 _07543_ (.A(_02765_),
    .B(_02767_),
    .Y(_02769_));
 sky130_fd_sc_hd__nor2_1 _07544_ (.A(_02768_),
    .B(_02769_),
    .Y(\u_decod.rs2_data_nxt[22] ));
 sky130_fd_sc_hd__nor2_1 _07545_ (.A(_01368_),
    .B(_01369_),
    .Y(_02770_));
 sky130_fd_sc_hd__or3b_1 _07546_ (.A(_01398_),
    .B(_02770_),
    .C_N(_02738_),
    .X(_02771_));
 sky130_fd_sc_hd__a21o_1 _07547_ (.A1(_01373_),
    .A2(_02738_),
    .B1(_01370_),
    .X(_02772_));
 sky130_fd_sc_hd__and4_1 _07548_ (.A(\u_decod.pc_q_o[21] ),
    .B(\u_decod.pc_q_o[22] ),
    .C(\u_decod.pc_q_o[23] ),
    .D(_02638_),
    .X(_02773_));
 sky130_fd_sc_hd__a31o_1 _07549_ (.A1(\u_decod.pc_q_o[21] ),
    .A2(\u_decod.pc_q_o[22] ),
    .A3(_02638_),
    .B1(\u_decod.pc_q_o[23] ),
    .X(_02774_));
 sky130_fd_sc_hd__and3b_1 _07550_ (.A_N(_02773_),
    .B(_01485_),
    .C(_02774_),
    .X(_02775_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_02619_),
    .B(net48),
    .Y(_02776_));
 sky130_fd_sc_hd__a21oi_1 _07552_ (.A1(_02618_),
    .A2(_02776_),
    .B1(_02621_),
    .Y(_02777_));
 sky130_fd_sc_hd__mux4_1 _07553_ (.A0(_01367_),
    .A1(_01289_),
    .A2(\u_decod.rs1_data_q[7] ),
    .A3(_01747_),
    .S0(_01468_),
    .S1(_01466_),
    .X(_02778_));
 sky130_fd_sc_hd__mux4_1 _07554_ (.A0(_02498_),
    .A1(_02584_),
    .A2(_02684_),
    .A3(_02778_),
    .S0(_01476_),
    .S1(_02685_),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _07555_ (.A0(_02734_),
    .A1(_02779_),
    .S(_02189_),
    .X(_02780_));
 sky130_fd_sc_hd__clkbuf_4 _07556_ (.A(\u_decod.instr_operation_q[1] ),
    .X(_02781_));
 sky130_fd_sc_hd__nor2_1 _07557_ (.A(_01368_),
    .B(_01820_),
    .Y(_02782_));
 sky130_fd_sc_hd__a221o_1 _07558_ (.A1(_02781_),
    .A2(_01369_),
    .B1(_02770_),
    .B2(_01435_),
    .C1(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__a22o_1 _07559_ (.A1(_01746_),
    .A2(_02780_),
    .B1(_02783_),
    .B2(_01260_),
    .X(_02784_));
 sky130_fd_sc_hd__o21a_1 _07560_ (.A1(_01467_),
    .A2(_02404_),
    .B1(_01498_),
    .X(_02785_));
 sky130_fd_sc_hd__mux2_1 _07561_ (.A0(_02579_),
    .A1(_02785_),
    .S(_01464_),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_1 _07562_ (.A0(_02680_),
    .A1(_02786_),
    .S(_02681_),
    .X(_02787_));
 sky130_fd_sc_hd__nor2_1 _07563_ (.A(_01480_),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__o211ai_2 _07564_ (.A1(_02781_),
    .A2(_01430_),
    .B1(\u_decod.instr_unit_q[1] ),
    .C1(_01427_),
    .Y(_02789_));
 sky130_fd_sc_hd__a211o_1 _07565_ (.A1(_01481_),
    .A2(_02728_),
    .B1(_02788_),
    .C1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__or4b_1 _07566_ (.A(_02775_),
    .B(_02777_),
    .C(_02784_),
    .D_N(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__a31o_2 _07567_ (.A1(_02332_),
    .A2(_02771_),
    .A3(_02772_),
    .B1(_02791_),
    .X(\u_decod.exe_ff_res_data_i[23] ));
 sky130_fd_sc_hd__a21o_1 _07568_ (.A1(\u_decod.dec0.instr_i[23] ),
    .A2(_01206_),
    .B1(_02646_),
    .X(_02792_));
 sky130_fd_sc_hd__a22o_1 _07569_ (.A1(\u_rf.reg30_q[23] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[23] ),
    .X(_02793_));
 sky130_fd_sc_hd__a221o_1 _07570_ (.A1(\u_rf.reg31_q[23] ),
    .A2(_01777_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[23] ),
    .C1(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__a22o_1 _07571_ (.A1(\u_rf.reg12_q[23] ),
    .A2(_01609_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[23] ),
    .X(_02795_));
 sky130_fd_sc_hd__a221o_1 _07572_ (.A1(\u_rf.reg9_q[23] ),
    .A2(_02360_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[23] ),
    .C1(_02795_),
    .X(_02796_));
 sky130_fd_sc_hd__a22o_1 _07573_ (.A1(\u_rf.reg6_q[23] ),
    .A2(_01557_),
    .B1(_01653_),
    .B2(\u_rf.reg22_q[23] ),
    .X(_02797_));
 sky130_fd_sc_hd__a221o_1 _07574_ (.A1(\u_rf.reg11_q[23] ),
    .A2(_02375_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[23] ),
    .C1(_02797_),
    .X(_02798_));
 sky130_fd_sc_hd__a22o_1 _07575_ (.A1(\u_rf.reg23_q[23] ),
    .A2(_02652_),
    .B1(_01791_),
    .B2(\u_rf.reg10_q[23] ),
    .X(_02799_));
 sky130_fd_sc_hd__a221o_1 _07576_ (.A1(\u_rf.reg13_q[23] ),
    .A2(_02376_),
    .B1(_01787_),
    .B2(\u_rf.reg18_q[23] ),
    .C1(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__or3_1 _07577_ (.A(_02796_),
    .B(_02798_),
    .C(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__a22o_1 _07578_ (.A1(\u_rf.reg16_q[23] ),
    .A2(_01565_),
    .B1(_01631_),
    .B2(\u_rf.reg17_q[23] ),
    .X(_02802_));
 sky130_fd_sc_hd__a221o_1 _07579_ (.A1(\u_rf.reg5_q[23] ),
    .A2(_02664_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[23] ),
    .C1(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__a22o_1 _07580_ (.A1(\u_rf.reg7_q[23] ),
    .A2(_01561_),
    .B1(_01606_),
    .B2(\u_rf.reg3_q[23] ),
    .X(_02804_));
 sky130_fd_sc_hd__a221o_1 _07581_ (.A1(\u_rf.reg0_q[23] ),
    .A2(_01664_),
    .B1(_02371_),
    .B2(\u_rf.reg15_q[23] ),
    .C1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__a22o_1 _07582_ (.A1(\u_rf.reg26_q[23] ),
    .A2(_02368_),
    .B1(_01645_),
    .B2(\u_rf.reg20_q[23] ),
    .X(_02806_));
 sky130_fd_sc_hd__a221o_1 _07583_ (.A1(\u_rf.reg25_q[23] ),
    .A2(_01783_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[23] ),
    .C1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__a22o_1 _07584_ (.A1(\u_rf.reg1_q[23] ),
    .A2(_02604_),
    .B1(_01659_),
    .B2(\u_rf.reg14_q[23] ),
    .X(_02808_));
 sky130_fd_sc_hd__a221o_1 _07585_ (.A1(\u_rf.reg29_q[23] ),
    .A2(_01780_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[23] ),
    .C1(_02808_),
    .X(_02809_));
 sky130_fd_sc_hd__or4_1 _07586_ (.A(_02803_),
    .B(_02805_),
    .C(_02807_),
    .D(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__o31a_2 _07587_ (.A1(_02794_),
    .A2(_02801_),
    .A3(_02810_),
    .B1(_02359_),
    .X(_02811_));
 sky130_fd_sc_hd__a221o_1 _07588_ (.A1(\u_decod.rf_ff_res_data_i[23] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_02792_),
    .C1(_02811_),
    .X(_02812_));
 sky130_fd_sc_hd__a21oi_1 _07589_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[23] ),
    .B1(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__nor2_1 _07590_ (.A(net200),
    .B(_02768_),
    .Y(_02814_));
 sky130_fd_sc_hd__xnor2_1 _07591_ (.A(_02813_),
    .B(_02814_),
    .Y(\u_decod.rs2_data_nxt[23] ));
 sky130_fd_sc_hd__nor2_1 _07592_ (.A(\u_decod.pc_q_o[24] ),
    .B(_02773_),
    .Y(_02815_));
 sky130_fd_sc_hd__and2_1 _07593_ (.A(\u_decod.pc_q_o[24] ),
    .B(_02773_),
    .X(_02816_));
 sky130_fd_sc_hd__a211o_1 _07594_ (.A1(_01372_),
    .A2(_01397_),
    .B1(_01369_),
    .C1(_01398_),
    .X(_02817_));
 sky130_fd_sc_hd__or2b_1 _07595_ (.A(_01368_),
    .B_N(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__and2_1 _07596_ (.A(_02818_),
    .B(_01405_),
    .X(_02819_));
 sky130_fd_sc_hd__inv_2 _07597_ (.A(_01280_),
    .Y(_02820_));
 sky130_fd_sc_hd__a221o_1 _07598_ (.A1(_02818_),
    .A2(_01375_),
    .B1(_02635_),
    .B2(_02819_),
    .C1(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__a211o_1 _07599_ (.A1(_01357_),
    .A2(_01393_),
    .B1(_01407_),
    .C1(_01280_),
    .X(_02822_));
 sky130_fd_sc_hd__and3_1 _07600_ (.A(\u_decod.rs2_data_q[24] ),
    .B(\u_decod.rs1_data_q[24] ),
    .C(_02781_),
    .X(_02823_));
 sky130_fd_sc_hd__a211o_1 _07601_ (.A1(_01278_),
    .A2(_01435_),
    .B1(_02823_),
    .C1(_01432_),
    .X(_02824_));
 sky130_fd_sc_hd__a32o_1 _07602_ (.A1(_01437_),
    .A2(_02821_),
    .A3(_02822_),
    .B1(_02824_),
    .B2(_01279_),
    .X(_02825_));
 sky130_fd_sc_hd__or2_1 _07603_ (.A(_01425_),
    .B(_02787_),
    .X(_02826_));
 sky130_fd_sc_hd__and3_1 _07604_ (.A(_01267_),
    .B(_01498_),
    .C(_02136_),
    .X(_02827_));
 sky130_fd_sc_hd__mux2_1 _07605_ (.A0(_02623_),
    .A1(_02827_),
    .S(_01472_),
    .X(_02828_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(_02681_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__o21a_1 _07607_ (.A1(_02681_),
    .A2(_02727_),
    .B1(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__nand2_1 _07608_ (.A(_02723_),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21bo_1 _07609_ (.A1(net49),
    .A2(net100),
    .B1_N(_02446_),
    .X(_02832_));
 sky130_fd_sc_hd__mux4_1 _07610_ (.A0(\u_decod.rs1_data_q[24] ),
    .A1(_01388_),
    .A2(\u_decod.rs1_data_q[8] ),
    .A3(_01061_),
    .S0(_01467_),
    .S1(_01461_),
    .X(_02833_));
 sky130_fd_sc_hd__mux2_1 _07611_ (.A0(_02629_),
    .A1(_02833_),
    .S(_01905_),
    .X(_02834_));
 sky130_fd_sc_hd__mux2_1 _07612_ (.A0(_02733_),
    .A1(_02834_),
    .S(_01476_),
    .X(_02835_));
 sky130_fd_sc_hd__mux2_1 _07613_ (.A0(_02779_),
    .A1(_02835_),
    .S(_01480_),
    .X(_02836_));
 sky130_fd_sc_hd__a22o_1 _07614_ (.A1(net133),
    .A2(_02832_),
    .B1(_02836_),
    .B2(_01746_),
    .X(_02837_));
 sky130_fd_sc_hd__a31o_1 _07615_ (.A1(_01443_),
    .A2(_02826_),
    .A3(_02831_),
    .B1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__a21oi_1 _07616_ (.A1(_01260_),
    .A2(_02825_),
    .B1(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__o31a_2 _07617_ (.A1(_02334_),
    .A2(_02815_),
    .A3(_02816_),
    .B1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__inv_2 _07618_ (.A(_02840_),
    .Y(\u_decod.exe_ff_res_data_i[24] ));
 sky130_fd_sc_hd__a21o_1 _07619_ (.A1(_01572_),
    .A2(_01224_),
    .B1(_02646_),
    .X(_02841_));
 sky130_fd_sc_hd__a22o_1 _07620_ (.A1(\u_rf.reg26_q[24] ),
    .A2(_02368_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[24] ),
    .X(_02842_));
 sky130_fd_sc_hd__a221o_1 _07621_ (.A1(\u_rf.reg24_q[24] ),
    .A2(_01784_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[24] ),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__a22o_1 _07622_ (.A1(\u_rf.reg30_q[24] ),
    .A2(_01581_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[24] ),
    .X(_02844_));
 sky130_fd_sc_hd__a221o_1 _07623_ (.A1(\u_rf.reg6_q[24] ),
    .A2(_01557_),
    .B1(_02376_),
    .B2(\u_rf.reg13_q[24] ),
    .C1(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__a22o_1 _07624_ (.A1(\u_rf.reg22_q[24] ),
    .A2(_01654_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[24] ),
    .X(_02846_));
 sky130_fd_sc_hd__a221o_1 _07625_ (.A1(\u_rf.reg11_q[24] ),
    .A2(_02375_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[24] ),
    .C1(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__a22o_1 _07626_ (.A1(\u_rf.reg25_q[24] ),
    .A2(_01783_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[24] ),
    .X(_02848_));
 sky130_fd_sc_hd__a221o_1 _07627_ (.A1(\u_rf.reg3_q[24] ),
    .A2(_02363_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[24] ),
    .C1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__or4_1 _07628_ (.A(_02843_),
    .B(_02845_),
    .C(_02847_),
    .D(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__a22o_1 _07629_ (.A1(\u_rf.reg21_q[24] ),
    .A2(_01639_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[24] ),
    .X(_02851_));
 sky130_fd_sc_hd__a221o_1 _07630_ (.A1(\u_rf.reg7_q[24] ),
    .A2(_01562_),
    .B1(_01780_),
    .B2(\u_rf.reg29_q[24] ),
    .C1(_02851_),
    .X(_02852_));
 sky130_fd_sc_hd__a22o_1 _07631_ (.A1(\u_rf.reg31_q[24] ),
    .A2(_01616_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[24] ),
    .X(_02853_));
 sky130_fd_sc_hd__a221o_1 _07632_ (.A1(\u_rf.reg0_q[24] ),
    .A2(_01664_),
    .B1(_01787_),
    .B2(\u_rf.reg18_q[24] ),
    .C1(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__a22o_1 _07633_ (.A1(\u_rf.reg16_q[24] ),
    .A2(_02307_),
    .B1(_01610_),
    .B2(\u_rf.reg12_q[24] ),
    .X(_02855_));
 sky130_fd_sc_hd__a221o_1 _07634_ (.A1(\u_rf.reg1_q[24] ),
    .A2(_02604_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[24] ),
    .C1(_02855_),
    .X(_02856_));
 sky130_fd_sc_hd__a22o_1 _07635_ (.A1(\u_rf.reg15_q[24] ),
    .A2(_02371_),
    .B1(_02652_),
    .B2(\u_rf.reg23_q[24] ),
    .X(_02857_));
 sky130_fd_sc_hd__a221o_1 _07636_ (.A1(\u_rf.reg5_q[24] ),
    .A2(_02664_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[24] ),
    .C1(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__or4_1 _07637_ (.A(_02852_),
    .B(_02854_),
    .C(_02856_),
    .D(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__o21a_1 _07638_ (.A1(_02850_),
    .A2(_02859_),
    .B1(_02359_),
    .X(_02860_));
 sky130_fd_sc_hd__a221oi_2 _07639_ (.A1(\u_decod.rf_ff_res_data_i[24] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_02841_),
    .C1(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__o21a_1 _07640_ (.A1(_01528_),
    .A2(_02840_),
    .B1(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__and4_1 _07641_ (.A(_02672_),
    .B(_02765_),
    .C(_02766_),
    .D(_02813_),
    .X(_02863_));
 sky130_fd_sc_hd__and3_1 _07642_ (.A(_02089_),
    .B(_02487_),
    .C(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__nor2_1 _07643_ (.A(net199),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__xnor2_1 _07644_ (.A(_02862_),
    .B(_02865_),
    .Y(\u_decod.rs2_data_nxt[24] ));
 sky130_fd_sc_hd__a21bo_1 _07645_ (.A1(_01278_),
    .A2(_02821_),
    .B1_N(_01277_),
    .X(_02866_));
 sky130_fd_sc_hd__nand3b_1 _07646_ (.A_N(_01277_),
    .B(_01278_),
    .C(_02821_),
    .Y(_02867_));
 sky130_fd_sc_hd__and3_1 _07647_ (.A(\u_decod.pc_q_o[24] ),
    .B(\u_decod.pc_q_o[25] ),
    .C(_02773_),
    .X(_02868_));
 sky130_fd_sc_hd__o21ai_1 _07648_ (.A1(\u_decod.pc_q_o[25] ),
    .A2(_02816_),
    .B1(_01485_),
    .Y(_02869_));
 sky130_fd_sc_hd__inv_2 _07649_ (.A(_02786_),
    .Y(_02870_));
 sky130_fd_sc_hd__o21ai_1 _07650_ (.A1(_01472_),
    .A2(_02679_),
    .B1(_01500_),
    .Y(_02871_));
 sky130_fd_sc_hd__mux2_1 _07651_ (.A0(_02870_),
    .A1(_02871_),
    .S(_02681_),
    .X(_02872_));
 sky130_fd_sc_hd__mux2_1 _07652_ (.A0(_02830_),
    .A1(_02872_),
    .S(_01425_),
    .X(_02873_));
 sky130_fd_sc_hd__mux4_1 _07653_ (.A0(\u_decod.rs1_data_q[25] ),
    .A1(_01380_),
    .A2(\u_decod.rs1_data_q[9] ),
    .A3(\u_decod.rs1_data_q[1] ),
    .S0(_01468_),
    .S1(_01466_),
    .X(_02874_));
 sky130_fd_sc_hd__mux4_1 _07654_ (.A0(_02584_),
    .A1(_02684_),
    .A2(_02778_),
    .A3(_02874_),
    .S0(_01475_),
    .S1(_02685_),
    .X(_02875_));
 sky130_fd_sc_hd__mux2_1 _07655_ (.A0(_02835_),
    .A1(_02875_),
    .S(_02189_),
    .X(_02876_));
 sky130_fd_sc_hd__and3_1 _07656_ (.A(\u_decod.rs2_data_q[25] ),
    .B(\u_decod.rs1_data_q[25] ),
    .C(_02781_),
    .X(_02877_));
 sky130_fd_sc_hd__a221o_1 _07657_ (.A1(_01430_),
    .A2(_01275_),
    .B1(_01277_),
    .B2(\u_decod.instr_operation_q[3] ),
    .C1(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__a22oi_1 _07658_ (.A1(_01506_),
    .A2(_02876_),
    .B1(_02878_),
    .B2(_01260_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _07659_ (.A(net100),
    .B(net50),
    .Y(_02880_));
 sky130_fd_sc_hd__a21o_1 _07660_ (.A1(_02618_),
    .A2(_02880_),
    .B1(_01057_),
    .X(_02881_));
 sky130_fd_sc_hd__o211a_1 _07661_ (.A1(_02789_),
    .A2(_02873_),
    .B1(_02879_),
    .C1(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__o21ai_1 _07662_ (.A1(_02868_),
    .A2(_02869_),
    .B1(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__a31o_1 _07663_ (.A1(_02332_),
    .A2(_02866_),
    .A3(_02867_),
    .B1(_02883_),
    .X(\u_decod.exe_ff_res_data_i[25] ));
 sky130_fd_sc_hd__a21o_1 _07664_ (.A1(\u_decod.dec0.funct7[0] ),
    .A2(_01206_),
    .B1(_02646_),
    .X(_02884_));
 sky130_fd_sc_hd__a22o_1 _07665_ (.A1(\u_rf.reg13_q[25] ),
    .A2(_01597_),
    .B1(_01656_),
    .B2(\u_rf.reg10_q[25] ),
    .X(_02885_));
 sky130_fd_sc_hd__a221o_1 _07666_ (.A1(\u_rf.reg6_q[25] ),
    .A2(_01556_),
    .B1(_01630_),
    .B2(\u_rf.reg17_q[25] ),
    .C1(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__a22o_1 _07667_ (.A1(\u_rf.reg7_q[25] ),
    .A2(_01560_),
    .B1(_01644_),
    .B2(\u_rf.reg20_q[25] ),
    .X(_02887_));
 sky130_fd_sc_hd__a221o_1 _07668_ (.A1(\u_rf.reg1_q[25] ),
    .A2(_01586_),
    .B1(_01671_),
    .B2(\u_rf.reg27_q[25] ),
    .C1(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__a22o_1 _07669_ (.A1(\u_rf.reg26_q[25] ),
    .A2(_01641_),
    .B1(_01649_),
    .B2(\u_rf.reg4_q[25] ),
    .X(_02889_));
 sky130_fd_sc_hd__a221o_1 _07670_ (.A1(\u_rf.reg12_q[25] ),
    .A2(_01609_),
    .B1(_01628_),
    .B2(\u_rf.reg29_q[25] ),
    .C1(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__a22o_1 _07671_ (.A1(\u_rf.reg15_q[25] ),
    .A2(_01600_),
    .B1(_01612_),
    .B2(\u_rf.reg23_q[25] ),
    .X(_02891_));
 sky130_fd_sc_hd__a221o_1 _07672_ (.A1(\u_rf.reg5_q[25] ),
    .A2(_01569_),
    .B1(_01606_),
    .B2(\u_rf.reg3_q[25] ),
    .C1(_02891_),
    .X(_02892_));
 sky130_fd_sc_hd__or4_1 _07673_ (.A(_02886_),
    .B(_02888_),
    .C(_02890_),
    .D(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__a22o_1 _07674_ (.A1(\u_rf.reg22_q[25] ),
    .A2(_01652_),
    .B1(_01673_),
    .B2(\u_rf.reg2_q[25] ),
    .X(_02894_));
 sky130_fd_sc_hd__a221o_1 _07675_ (.A1(\u_rf.reg31_q[25] ),
    .A2(_01616_),
    .B1(_01658_),
    .B2(\u_rf.reg14_q[25] ),
    .C1(_02894_),
    .X(_02895_));
 sky130_fd_sc_hd__a22o_1 _07676_ (.A1(\u_rf.reg25_q[25] ),
    .A2(_01575_),
    .B1(_01621_),
    .B2(\u_rf.reg24_q[25] ),
    .X(_02896_));
 sky130_fd_sc_hd__a221o_1 _07677_ (.A1(\u_rf.reg18_q[25] ),
    .A2(_01592_),
    .B1(_01638_),
    .B2(\u_rf.reg21_q[25] ),
    .C1(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__a22o_1 _07678_ (.A1(\u_rf.reg0_q[25] ),
    .A2(_01662_),
    .B1(_01666_),
    .B2(\u_rf.reg8_q[25] ),
    .X(_02898_));
 sky130_fd_sc_hd__a221o_1 _07679_ (.A1(\u_rf.reg16_q[25] ),
    .A2(_01564_),
    .B1(_01636_),
    .B2(\u_rf.reg9_q[25] ),
    .C1(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__a22o_1 _07680_ (.A1(\u_rf.reg30_q[25] ),
    .A2(_01579_),
    .B1(_01624_),
    .B2(\u_rf.reg28_q[25] ),
    .X(_02900_));
 sky130_fd_sc_hd__a221o_1 _07681_ (.A1(\u_rf.reg11_q[25] ),
    .A2(_01584_),
    .B1(_01595_),
    .B2(\u_rf.reg19_q[25] ),
    .C1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__or4_1 _07682_ (.A(_02895_),
    .B(_02897_),
    .C(_02899_),
    .D(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__or2_1 _07683_ (.A(_02893_),
    .B(_02902_),
    .X(_02903_));
 sky130_fd_sc_hd__and2_1 _07684_ (.A(_01680_),
    .B(_02903_),
    .X(_02904_));
 sky130_fd_sc_hd__a221o_1 _07685_ (.A1(\u_decod.rf_ff_res_data_i[25] ),
    .A2(_01550_),
    .B1(_02743_),
    .B2(_02884_),
    .C1(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__a21oi_1 _07686_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[25] ),
    .B1(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__a21oi_1 _07687_ (.A1(_02862_),
    .A2(_02864_),
    .B1(net200),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_1 _07688_ (.A(_02906_),
    .B(_02907_),
    .Y(\u_decod.rs2_data_nxt[25] ));
 sky130_fd_sc_hd__nor2_1 _07689_ (.A(\u_decod.pc_q_o[26] ),
    .B(_02868_),
    .Y(_02908_));
 sky130_fd_sc_hd__and2_1 _07690_ (.A(\u_decod.pc_q_o[26] ),
    .B(_02868_),
    .X(_02909_));
 sky130_fd_sc_hd__inv_2 _07691_ (.A(_01286_),
    .Y(_02910_));
 sky130_fd_sc_hd__a311o_1 _07692_ (.A1(_01276_),
    .A2(_01278_),
    .A3(_02821_),
    .B1(_02910_),
    .C1(_01410_),
    .X(_02911_));
 sky130_fd_sc_hd__a21o_1 _07693_ (.A1(_01357_),
    .A2(_01393_),
    .B1(_01407_),
    .X(_02912_));
 sky130_fd_sc_hd__a311o_1 _07694_ (.A1(_01277_),
    .A2(_01280_),
    .A3(_02912_),
    .B1(_01411_),
    .C1(_01286_),
    .X(_02913_));
 sky130_fd_sc_hd__a21o_1 _07695_ (.A1(_01285_),
    .A2(_01435_),
    .B1(_01432_),
    .X(_02914_));
 sky130_fd_sc_hd__a22o_1 _07696_ (.A1(_02781_),
    .A2(_01409_),
    .B1(_02914_),
    .B2(_01284_),
    .X(_02915_));
 sky130_fd_sc_hd__a31o_1 _07697_ (.A1(_02332_),
    .A2(_02911_),
    .A3(_02913_),
    .B1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__mux4_1 _07698_ (.A0(\u_decod.rs1_data_q[26] ),
    .A1(_01384_),
    .A2(_01302_),
    .A3(\u_decod.rs1_data_q[2] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _07699_ (.A0(_02732_),
    .A1(_02917_),
    .S(_02685_),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _07700_ (.A0(_02834_),
    .A1(_02918_),
    .S(_01477_),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _07701_ (.A0(_02875_),
    .A1(_02919_),
    .S(_01481_),
    .X(_02920_));
 sky130_fd_sc_hd__o21a_1 _07702_ (.A1(_01472_),
    .A2(_02725_),
    .B1(_01500_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _07703_ (.A0(_02828_),
    .A1(_02921_),
    .S(_02681_),
    .X(_02922_));
 sky130_fd_sc_hd__o21ai_1 _07704_ (.A1(_01481_),
    .A2(_02922_),
    .B1(_01443_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21oi_1 _07705_ (.A1(_01481_),
    .A2(_02872_),
    .B1(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _07706_ (.A(_02619_),
    .B(net51),
    .Y(_02925_));
 sky130_fd_sc_hd__a21oi_1 _07707_ (.A1(_02618_),
    .A2(_02925_),
    .B1(_02621_),
    .Y(_02926_));
 sky130_fd_sc_hd__a211o_1 _07708_ (.A1(_01746_),
    .A2(_02920_),
    .B1(_02924_),
    .C1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__a21oi_1 _07709_ (.A1(_01260_),
    .A2(_02916_),
    .B1(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__o31a_2 _07710_ (.A1(_02334_),
    .A2(_02908_),
    .A3(_02909_),
    .B1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__inv_2 _07711_ (.A(_02929_),
    .Y(\u_decod.exe_ff_res_data_i[26] ));
 sky130_fd_sc_hd__a21o_1 _07712_ (.A1(\u_decod.dec0.funct7[1] ),
    .A2(_01224_),
    .B1(_02646_),
    .X(_02930_));
 sky130_fd_sc_hd__a22o_1 _07713_ (.A1(\u_rf.reg15_q[26] ),
    .A2(_01601_),
    .B1(_02363_),
    .B2(\u_rf.reg3_q[26] ),
    .X(_02931_));
 sky130_fd_sc_hd__a221o_1 _07714_ (.A1(\u_rf.reg7_q[26] ),
    .A2(_01562_),
    .B1(_02604_),
    .B2(\u_rf.reg1_q[26] ),
    .C1(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__a22o_1 _07715_ (.A1(\u_rf.reg13_q[26] ),
    .A2(_01598_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[26] ),
    .X(_02933_));
 sky130_fd_sc_hd__a221o_1 _07716_ (.A1(\u_rf.reg10_q[26] ),
    .A2(_02380_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[26] ),
    .C1(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__a22o_1 _07717_ (.A1(\u_rf.reg12_q[26] ),
    .A2(_01609_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[26] ),
    .X(_02935_));
 sky130_fd_sc_hd__a221o_1 _07718_ (.A1(\u_rf.reg29_q[26] ),
    .A2(_01780_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[26] ),
    .C1(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__a22o_1 _07719_ (.A1(\u_rf.reg6_q[26] ),
    .A2(_01557_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[26] ),
    .X(_02937_));
 sky130_fd_sc_hd__a221o_1 _07720_ (.A1(\u_rf.reg5_q[26] ),
    .A2(_02664_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[26] ),
    .C1(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__or4_1 _07721_ (.A(_02932_),
    .B(_02934_),
    .C(_02936_),
    .D(_02938_),
    .X(_02939_));
 sky130_fd_sc_hd__a22o_1 _07722_ (.A1(\u_rf.reg16_q[26] ),
    .A2(_01565_),
    .B1(_02652_),
    .B2(\u_rf.reg23_q[26] ),
    .X(_02940_));
 sky130_fd_sc_hd__a221o_1 _07723_ (.A1(\u_rf.reg17_q[26] ),
    .A2(_02379_),
    .B1(_02360_),
    .B2(\u_rf.reg9_q[26] ),
    .C1(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__a22o_1 _07724_ (.A1(\u_rf.reg30_q[26] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[26] ),
    .X(_02942_));
 sky130_fd_sc_hd__a221o_1 _07725_ (.A1(\u_rf.reg22_q[26] ),
    .A2(_01654_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[26] ),
    .C1(_02942_),
    .X(_02943_));
 sky130_fd_sc_hd__a22o_1 _07726_ (.A1(\u_rf.reg0_q[26] ),
    .A2(_01663_),
    .B1(_01674_),
    .B2(\u_rf.reg2_q[26] ),
    .X(_02944_));
 sky130_fd_sc_hd__a221o_1 _07727_ (.A1(\u_rf.reg31_q[26] ),
    .A2(_01777_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[26] ),
    .C1(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__a22o_1 _07728_ (.A1(\u_rf.reg18_q[26] ),
    .A2(_01787_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[26] ),
    .X(_02946_));
 sky130_fd_sc_hd__a221o_1 _07729_ (.A1(\u_rf.reg25_q[26] ),
    .A2(_01783_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[26] ),
    .C1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__or4_1 _07730_ (.A(_02941_),
    .B(_02943_),
    .C(_02945_),
    .D(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__or2_1 _07731_ (.A(_02939_),
    .B(_02948_),
    .X(_02949_));
 sky130_fd_sc_hd__and2_1 _07732_ (.A(_02359_),
    .B(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__a221oi_2 _07733_ (.A1(\u_decod.rf_ff_res_data_i[26] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_02930_),
    .C1(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__o21a_1 _07734_ (.A1(_01528_),
    .A2(_02929_),
    .B1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__o211a_1 _07735_ (.A1(_01528_),
    .A2(_02840_),
    .B1(_02861_),
    .C1(_02906_),
    .X(_02953_));
 sky130_fd_sc_hd__a21oi_1 _07736_ (.A1(_02864_),
    .A2(_02953_),
    .B1(net200),
    .Y(_02954_));
 sky130_fd_sc_hd__xnor2_1 _07737_ (.A(_02952_),
    .B(_02954_),
    .Y(\u_decod.rs2_data_nxt[26] ));
 sky130_fd_sc_hd__a21bo_1 _07738_ (.A1(_01285_),
    .A2(_02911_),
    .B1_N(_01283_),
    .X(_02955_));
 sky130_fd_sc_hd__or3b_1 _07739_ (.A(_01283_),
    .B(_01409_),
    .C_N(_02911_),
    .X(_02956_));
 sky130_fd_sc_hd__or2_1 _07740_ (.A(\u_decod.pc_q_o[27] ),
    .B(_02909_),
    .X(_02957_));
 sky130_fd_sc_hd__nand2_1 _07741_ (.A(\u_decod.pc_q_o[27] ),
    .B(_02909_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21bo_1 _07742_ (.A1(_02619_),
    .A2(net52),
    .B1_N(_02618_),
    .X(_02959_));
 sky130_fd_sc_hd__o21ai_1 _07743_ (.A1(_01472_),
    .A2(_02785_),
    .B1(_01500_),
    .Y(_02960_));
 sky130_fd_sc_hd__mux2_1 _07744_ (.A0(_02871_),
    .A1(_02960_),
    .S(_02681_),
    .X(_02961_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_02723_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__o211a_1 _07746_ (.A1(_02723_),
    .A2(_02922_),
    .B1(_02962_),
    .C1(_01443_),
    .X(_02963_));
 sky130_fd_sc_hd__mux4_1 _07747_ (.A0(\u_decod.rs1_data_q[27] ),
    .A1(_01376_),
    .A2(\u_decod.rs1_data_q[11] ),
    .A3(\u_decod.rs1_data_q[3] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_02964_));
 sky130_fd_sc_hd__mux4_1 _07748_ (.A0(_02684_),
    .A1(_02778_),
    .A2(_02874_),
    .A3(_02964_),
    .S0(_01476_),
    .S1(_02685_),
    .X(_02965_));
 sky130_fd_sc_hd__mux2_1 _07749_ (.A0(_02919_),
    .A1(_02965_),
    .S(_01481_),
    .X(_02966_));
 sky130_fd_sc_hd__and3_1 _07750_ (.A(\u_decod.rs2_data_q[27] ),
    .B(\u_decod.rs1_data_q[27] ),
    .C(_02781_),
    .X(_02967_));
 sky130_fd_sc_hd__a221o_1 _07751_ (.A1(_01430_),
    .A2(_01282_),
    .B1(_01283_),
    .B2(\u_decod.instr_operation_q[3] ),
    .C1(_02967_),
    .X(_02968_));
 sky130_fd_sc_hd__a22o_1 _07752_ (.A1(_01746_),
    .A2(_02966_),
    .B1(_02968_),
    .B2(_01260_),
    .X(_02969_));
 sky130_fd_sc_hd__a211o_1 _07753_ (.A1(net133),
    .A2(_02959_),
    .B1(_02963_),
    .C1(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__a31o_1 _07754_ (.A1(_01485_),
    .A2(_02957_),
    .A3(_02958_),
    .B1(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__a31oi_2 _07755_ (.A1(_02332_),
    .A2(_02955_),
    .A3(_02956_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__inv_2 _07756_ (.A(_02972_),
    .Y(\u_decod.exe_ff_res_data_i[27] ));
 sky130_fd_sc_hd__a21o_1 _07757_ (.A1(\u_decod.dec0.funct7[2] ),
    .A2(_01224_),
    .B1(_02646_),
    .X(_02973_));
 sky130_fd_sc_hd__a22o_1 _07758_ (.A1(\u_rf.reg27_q[27] ),
    .A2(_02386_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[27] ),
    .X(_02974_));
 sky130_fd_sc_hd__a221o_1 _07759_ (.A1(\u_rf.reg13_q[27] ),
    .A2(_02376_),
    .B1(_01787_),
    .B2(\u_rf.reg18_q[27] ),
    .C1(_02974_),
    .X(_02975_));
 sky130_fd_sc_hd__a22o_1 _07760_ (.A1(\u_rf.reg31_q[27] ),
    .A2(_01777_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[27] ),
    .X(_02976_));
 sky130_fd_sc_hd__a221o_1 _07761_ (.A1(\u_rf.reg12_q[27] ),
    .A2(_01610_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[27] ),
    .C1(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__a22o_1 _07762_ (.A1(\u_rf.reg6_q[27] ),
    .A2(_01557_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[27] ),
    .X(_02978_));
 sky130_fd_sc_hd__a221o_1 _07763_ (.A1(\u_rf.reg23_q[27] ),
    .A2(_02652_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[27] ),
    .C1(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__a22o_1 _07764_ (.A1(\u_rf.reg30_q[27] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[27] ),
    .X(_02980_));
 sky130_fd_sc_hd__a221o_1 _07765_ (.A1(\u_rf.reg9_q[27] ),
    .A2(_02360_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[27] ),
    .C1(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__or4_1 _07766_ (.A(_02975_),
    .B(_02977_),
    .C(_02979_),
    .D(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__a22o_1 _07767_ (.A1(\u_rf.reg16_q[27] ),
    .A2(_02307_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[27] ),
    .X(_02983_));
 sky130_fd_sc_hd__a221o_1 _07768_ (.A1(\u_rf.reg5_q[27] ),
    .A2(_02664_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[27] ),
    .C1(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__a22o_1 _07769_ (.A1(\u_rf.reg7_q[27] ),
    .A2(_01562_),
    .B1(_02363_),
    .B2(\u_rf.reg3_q[27] ),
    .X(_02985_));
 sky130_fd_sc_hd__a221o_1 _07770_ (.A1(\u_rf.reg0_q[27] ),
    .A2(_01664_),
    .B1(_02371_),
    .B2(\u_rf.reg15_q[27] ),
    .C1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__a22o_1 _07771_ (.A1(\u_rf.reg1_q[27] ),
    .A2(_02604_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[27] ),
    .X(_02987_));
 sky130_fd_sc_hd__a221o_1 _07772_ (.A1(\u_rf.reg29_q[27] ),
    .A2(_01780_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[27] ),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__a22o_1 _07773_ (.A1(\u_rf.reg26_q[27] ),
    .A2(_02368_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[27] ),
    .X(_02989_));
 sky130_fd_sc_hd__a221o_1 _07774_ (.A1(\u_rf.reg25_q[27] ),
    .A2(_01783_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[27] ),
    .C1(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__or4_1 _07775_ (.A(_02984_),
    .B(_02986_),
    .C(_02988_),
    .D(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o21a_1 _07776_ (.A1(_02982_),
    .A2(_02991_),
    .B1(_02359_),
    .X(_02992_));
 sky130_fd_sc_hd__a221o_1 _07777_ (.A1(\u_decod.rf_ff_res_data_i[27] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_02973_),
    .C1(_02992_),
    .X(_02993_));
 sky130_fd_sc_hd__a21oi_1 _07778_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[27] ),
    .B1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__o211a_1 _07779_ (.A1(_01528_),
    .A2(_02929_),
    .B1(_02951_),
    .C1(_02953_),
    .X(_02995_));
 sky130_fd_sc_hd__and4_1 _07780_ (.A(_02089_),
    .B(_02487_),
    .C(_02863_),
    .D(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__nor2_1 _07781_ (.A(_02229_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__xnor2_1 _07782_ (.A(_02994_),
    .B(_02997_),
    .Y(\u_decod.rs2_data_nxt[27] ));
 sky130_fd_sc_hd__a21oi_1 _07783_ (.A1(\u_decod.pc_q_o[27] ),
    .A2(_02909_),
    .B1(\u_decod.pc_q_o[28] ),
    .Y(_02998_));
 sky130_fd_sc_hd__and3_1 _07784_ (.A(\u_decod.pc_q_o[27] ),
    .B(\u_decod.pc_q_o[28] ),
    .C(_02909_),
    .X(_02999_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(_02781_),
    .B(_01264_),
    .Y(_03000_));
 sky130_fd_sc_hd__o211a_1 _07786_ (.A1(_01264_),
    .A2(_02244_),
    .B1(_03000_),
    .C1(_01820_),
    .X(_03001_));
 sky130_fd_sc_hd__a21oi_1 _07787_ (.A1(_01357_),
    .A2(_01393_),
    .B1(_01407_),
    .Y(_03002_));
 sky130_fd_sc_hd__o21ai_2 _07788_ (.A1(_01287_),
    .A2(_03002_),
    .B1(_01413_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _07789_ (.A(_01266_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__o21a_1 _07790_ (.A1(_01266_),
    .A2(_03003_),
    .B1(_02332_),
    .X(_03005_));
 sky130_fd_sc_hd__a2bb2o_1 _07791_ (.A1_N(_01265_),
    .A2_N(_03001_),
    .B1(_03004_),
    .B2(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__a21bo_1 _07792_ (.A1(_02619_),
    .A2(net53),
    .B1_N(_02618_),
    .X(_03007_));
 sky130_fd_sc_hd__inv_2 _07793_ (.A(_02961_),
    .Y(_03008_));
 sky130_fd_sc_hd__and2_1 _07794_ (.A(_01500_),
    .B(_02827_),
    .X(_03009_));
 sky130_fd_sc_hd__mux2_1 _07795_ (.A0(_02921_),
    .A1(_03009_),
    .S(_02681_),
    .X(_03010_));
 sky130_fd_sc_hd__mux2_1 _07796_ (.A0(_03008_),
    .A1(_03010_),
    .S(_02723_),
    .X(_03011_));
 sky130_fd_sc_hd__mux4_1 _07797_ (.A0(\u_decod.rs1_data_q[28] ),
    .A1(_01363_),
    .A2(_01297_),
    .A3(\u_decod.rs1_data_q[4] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_03012_));
 sky130_fd_sc_hd__mux2_1 _07798_ (.A0(_02833_),
    .A1(_03012_),
    .S(_02685_),
    .X(_03013_));
 sky130_fd_sc_hd__mux2_1 _07799_ (.A0(_02918_),
    .A1(_03013_),
    .S(_01477_),
    .X(_03014_));
 sky130_fd_sc_hd__mux2_1 _07800_ (.A0(_02965_),
    .A1(_03014_),
    .S(_01481_),
    .X(_03015_));
 sky130_fd_sc_hd__a22o_1 _07801_ (.A1(_01443_),
    .A2(_03011_),
    .B1(_03015_),
    .B2(_01746_),
    .X(_03016_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(net133),
    .A2(_03007_),
    .B1(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__a21oi_1 _07803_ (.A1(_01260_),
    .A2(_03006_),
    .B1(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__o31a_1 _07804_ (.A1(_02334_),
    .A2(_02998_),
    .A3(_02999_),
    .B1(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__inv_2 _07805_ (.A(_03019_),
    .Y(\u_decod.exe_ff_res_data_i[28] ));
 sky130_fd_sc_hd__a21o_1 _07806_ (.A1(\u_decod.dec0.funct7[3] ),
    .A2(_01224_),
    .B1(_02646_),
    .X(_03020_));
 sky130_fd_sc_hd__a22o_1 _07807_ (.A1(\u_rf.reg10_q[28] ),
    .A2(_02380_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[28] ),
    .X(_03021_));
 sky130_fd_sc_hd__a221o_1 _07808_ (.A1(\u_rf.reg21_q[28] ),
    .A2(_02364_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[28] ),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__a22o_1 _07809_ (.A1(\u_rf.reg25_q[28] ),
    .A2(_01783_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[28] ),
    .X(_03023_));
 sky130_fd_sc_hd__a221o_1 _07810_ (.A1(\u_rf.reg7_q[28] ),
    .A2(_01562_),
    .B1(_01780_),
    .B2(\u_rf.reg29_q[28] ),
    .C1(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__a22o_1 _07811_ (.A1(\u_rf.reg19_q[28] ),
    .A2(_02665_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[28] ),
    .X(_03025_));
 sky130_fd_sc_hd__a221o_1 _07812_ (.A1(\u_rf.reg12_q[28] ),
    .A2(_01610_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[28] ),
    .C1(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__a22o_1 _07813_ (.A1(\u_rf.reg30_q[28] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[28] ),
    .X(_03027_));
 sky130_fd_sc_hd__a221o_1 _07814_ (.A1(\u_rf.reg0_q[28] ),
    .A2(_01664_),
    .B1(_02371_),
    .B2(\u_rf.reg15_q[28] ),
    .C1(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__or4_1 _07815_ (.A(_03022_),
    .B(_03024_),
    .C(_03026_),
    .D(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__a22o_1 _07816_ (.A1(\u_rf.reg6_q[28] ),
    .A2(_01557_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[28] ),
    .X(_03030_));
 sky130_fd_sc_hd__a221o_1 _07817_ (.A1(\u_rf.reg23_q[28] ),
    .A2(_02652_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[28] ),
    .C1(_03030_),
    .X(_03031_));
 sky130_fd_sc_hd__a22o_1 _07818_ (.A1(\u_rf.reg5_q[28] ),
    .A2(_02664_),
    .B1(_02360_),
    .B2(\u_rf.reg9_q[28] ),
    .X(_03032_));
 sky130_fd_sc_hd__a221o_1 _07819_ (.A1(\u_rf.reg3_q[28] ),
    .A2(_02363_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[28] ),
    .C1(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__a22o_1 _07820_ (.A1(\u_rf.reg1_q[28] ),
    .A2(_02604_),
    .B1(_02376_),
    .B2(\u_rf.reg13_q[28] ),
    .X(_03034_));
 sky130_fd_sc_hd__a221o_1 _07821_ (.A1(\u_rf.reg31_q[28] ),
    .A2(_01777_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[28] ),
    .C1(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__a22o_1 _07822_ (.A1(\u_rf.reg16_q[28] ),
    .A2(_02307_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[28] ),
    .X(_03036_));
 sky130_fd_sc_hd__a221o_1 _07823_ (.A1(\u_rf.reg18_q[28] ),
    .A2(_01787_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[28] ),
    .C1(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__or4_1 _07824_ (.A(_03031_),
    .B(_03033_),
    .C(_03035_),
    .D(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__o21a_1 _07825_ (.A1(_03029_),
    .A2(_03038_),
    .B1(_02359_),
    .X(_03039_));
 sky130_fd_sc_hd__a221o_1 _07826_ (.A1(\u_decod.rf_ff_res_data_i[28] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_03020_),
    .C1(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__a21o_1 _07827_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[28] ),
    .B1(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_02994_),
    .B(_02996_),
    .Y(_03042_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(_01897_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor2_1 _07830_ (.A(_03041_),
    .B(_03043_),
    .Y(\u_decod.rs2_data_nxt[28] ));
 sky130_fd_sc_hd__a21oi_1 _07831_ (.A1(_01266_),
    .A2(_03003_),
    .B1(_01264_),
    .Y(_03044_));
 sky130_fd_sc_hd__xnor2_1 _07832_ (.A(_01263_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__and3_1 _07833_ (.A(\u_decod.rs2_data_q[29] ),
    .B(\u_decod.rs1_data_q[29] ),
    .C(_02781_),
    .X(_03046_));
 sky130_fd_sc_hd__a221o_1 _07834_ (.A1(\u_decod.instr_operation_q[3] ),
    .A2(_01263_),
    .B1(_01432_),
    .B2(_01414_),
    .C1(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__a21boi_1 _07835_ (.A1(_01477_),
    .A2(_02960_),
    .B1_N(_01502_),
    .Y(_03048_));
 sky130_fd_sc_hd__mux2_1 _07836_ (.A0(_03010_),
    .A1(_03048_),
    .S(_02723_),
    .X(_03049_));
 sky130_fd_sc_hd__a21bo_1 _07837_ (.A1(_02619_),
    .A2(net54),
    .B1_N(_02618_),
    .X(_03050_));
 sky130_fd_sc_hd__mux4_1 _07838_ (.A0(\u_decod.rs1_data_q[29] ),
    .A1(_01358_),
    .A2(\u_decod.rs1_data_q[13] ),
    .A3(\u_decod.rs1_data_q[5] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_03051_));
 sky130_fd_sc_hd__mux4_1 _07839_ (.A0(_02778_),
    .A1(_02874_),
    .A2(_02964_),
    .A3(_03051_),
    .S0(_01477_),
    .S1(_02685_),
    .X(_03052_));
 sky130_fd_sc_hd__mux2_1 _07840_ (.A0(_03014_),
    .A1(_03052_),
    .S(_01481_),
    .X(_03053_));
 sky130_fd_sc_hd__a22o_1 _07841_ (.A1(net133),
    .A2(_03050_),
    .B1(_03053_),
    .B2(_01746_),
    .X(_03054_));
 sky130_fd_sc_hd__a21o_1 _07842_ (.A1(_01443_),
    .A2(_03049_),
    .B1(_03054_),
    .X(_03055_));
 sky130_fd_sc_hd__o21ai_1 _07843_ (.A1(\u_decod.pc_q_o[29] ),
    .A2(_02999_),
    .B1(_01485_),
    .Y(_03056_));
 sky130_fd_sc_hd__a21oi_1 _07844_ (.A1(\u_decod.pc_q_o[29] ),
    .A2(_02999_),
    .B1(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__a211o_1 _07845_ (.A1(_01260_),
    .A2(_03047_),
    .B1(_03055_),
    .C1(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__a21oi_1 _07846_ (.A1(_02332_),
    .A2(_03045_),
    .B1(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__inv_2 _07847_ (.A(_03059_),
    .Y(\u_decod.exe_ff_res_data_i[29] ));
 sky130_fd_sc_hd__a21o_1 _07848_ (.A1(\u_decod.dec0.funct7[4] ),
    .A2(_01224_),
    .B1(_02646_),
    .X(_03060_));
 sky130_fd_sc_hd__a22o_1 _07849_ (.A1(\u_rf.reg18_q[29] ),
    .A2(_01787_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[29] ),
    .X(_03061_));
 sky130_fd_sc_hd__a221o_1 _07850_ (.A1(\u_rf.reg13_q[29] ),
    .A2(_02376_),
    .B1(_01777_),
    .B2(\u_rf.reg31_q[29] ),
    .C1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__a22o_1 _07851_ (.A1(\u_rf.reg0_q[29] ),
    .A2(_01664_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[29] ),
    .X(_03063_));
 sky130_fd_sc_hd__a221o_1 _07852_ (.A1(\u_rf.reg5_q[29] ),
    .A2(_02664_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[29] ),
    .C1(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__a22o_1 _07853_ (.A1(\u_rf.reg24_q[29] ),
    .A2(_01784_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[29] ),
    .X(_03065_));
 sky130_fd_sc_hd__a221o_1 _07854_ (.A1(\u_rf.reg25_q[29] ),
    .A2(_01783_),
    .B1(_02652_),
    .B2(\u_rf.reg23_q[29] ),
    .C1(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__a22o_1 _07855_ (.A1(\u_rf.reg7_q[29] ),
    .A2(_01562_),
    .B1(_02363_),
    .B2(\u_rf.reg3_q[29] ),
    .X(_03067_));
 sky130_fd_sc_hd__a221o_1 _07856_ (.A1(\u_rf.reg16_q[29] ),
    .A2(_02307_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[29] ),
    .C1(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__or4_1 _07857_ (.A(_03062_),
    .B(_03064_),
    .C(_03066_),
    .D(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__a22o_1 _07858_ (.A1(\u_rf.reg28_q[29] ),
    .A2(_02419_),
    .B1(_02360_),
    .B2(\u_rf.reg9_q[29] ),
    .X(_03070_));
 sky130_fd_sc_hd__a221o_1 _07859_ (.A1(\u_rf.reg29_q[29] ),
    .A2(_01780_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[29] ),
    .C1(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__a22o_1 _07860_ (.A1(\u_rf.reg1_q[29] ),
    .A2(_02604_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[29] ),
    .X(_03072_));
 sky130_fd_sc_hd__a221o_1 _07861_ (.A1(\u_rf.reg15_q[29] ),
    .A2(_02371_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[29] ),
    .C1(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__a22o_1 _07862_ (.A1(\u_rf.reg12_q[29] ),
    .A2(_01610_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[29] ),
    .X(_03074_));
 sky130_fd_sc_hd__a221o_1 _07863_ (.A1(\u_rf.reg11_q[29] ),
    .A2(_02375_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[29] ),
    .C1(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__a22o_1 _07864_ (.A1(\u_rf.reg6_q[29] ),
    .A2(_01557_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[29] ),
    .X(_03076_));
 sky130_fd_sc_hd__a221o_1 _07865_ (.A1(\u_rf.reg30_q[29] ),
    .A2(_01581_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[29] ),
    .C1(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__or4_1 _07866_ (.A(_03071_),
    .B(_03073_),
    .C(_03075_),
    .D(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__o21a_1 _07867_ (.A1(_03069_),
    .A2(_03078_),
    .B1(_02359_),
    .X(_03079_));
 sky130_fd_sc_hd__a221o_1 _07868_ (.A1(\u_decod.rf_ff_res_data_i[29] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_03060_),
    .C1(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__a21o_1 _07869_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[29] ),
    .B1(_03080_),
    .X(_03081_));
 sky130_fd_sc_hd__o21ai_1 _07870_ (.A1(_03041_),
    .A2(_03042_),
    .B1(_01897_),
    .Y(_03082_));
 sky130_fd_sc_hd__xnor2_1 _07871_ (.A(_03081_),
    .B(_03082_),
    .Y(\u_decod.rs2_data_nxt[29] ));
 sky130_fd_sc_hd__a31o_1 _07872_ (.A1(_01263_),
    .A2(_01266_),
    .A3(_03003_),
    .B1(_01415_),
    .X(_03083_));
 sky130_fd_sc_hd__nor2_1 _07873_ (.A(_01273_),
    .B(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__a21o_1 _07874_ (.A1(_01273_),
    .A2(_03083_),
    .B1(_01765_),
    .X(_03085_));
 sky130_fd_sc_hd__a21oi_1 _07875_ (.A1(\u_decod.pc_q_o[29] ),
    .A2(_02999_),
    .B1(\u_decod.pc_q_o[30] ),
    .Y(_03086_));
 sky130_fd_sc_hd__and3_1 _07876_ (.A(\u_decod.pc_q_o[29] ),
    .B(\u_decod.pc_q_o[30] ),
    .C(_02999_),
    .X(_03087_));
 sky130_fd_sc_hd__nand3_1 _07877_ (.A(\u_decod.instr_operation_q[0] ),
    .B(\u_decod.instr_unit_q[1] ),
    .C(_01427_),
    .Y(_03088_));
 sky130_fd_sc_hd__inv_2 _07878_ (.A(_03052_),
    .Y(_03089_));
 sky130_fd_sc_hd__mux4_1 _07879_ (.A0(\u_decod.rs1_data_q[30] ),
    .A1(_01371_),
    .A2(_01292_),
    .A3(\u_decod.rs1_data_q[6] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_03090_));
 sky130_fd_sc_hd__mux2_1 _07880_ (.A0(_02917_),
    .A1(_03090_),
    .S(_02685_),
    .X(_03091_));
 sky130_fd_sc_hd__or2_1 _07881_ (.A(_02681_),
    .B(_03091_),
    .X(_03092_));
 sky130_fd_sc_hd__o21ai_1 _07882_ (.A1(_01477_),
    .A2(_03013_),
    .B1(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__mux2_1 _07883_ (.A0(_03089_),
    .A1(_03093_),
    .S(_01481_),
    .X(_03094_));
 sky130_fd_sc_hd__o21a_1 _07884_ (.A1(_01272_),
    .A2(_02244_),
    .B1(_01820_),
    .X(_03095_));
 sky130_fd_sc_hd__o2bb2a_1 _07885_ (.A1_N(_01272_),
    .A2_N(_01429_),
    .B1(_03095_),
    .B2(_01271_),
    .X(_03096_));
 sky130_fd_sc_hd__nand2_1 _07886_ (.A(_02619_),
    .B(net56),
    .Y(_03097_));
 sky130_fd_sc_hd__a21o_1 _07887_ (.A1(_02618_),
    .A2(_03097_),
    .B1(_02621_),
    .X(_03098_));
 sky130_fd_sc_hd__nand2_1 _07888_ (.A(_01502_),
    .B(_03009_),
    .Y(_03099_));
 sky130_fd_sc_hd__nor2_1 _07889_ (.A(_02723_),
    .B(_03048_),
    .Y(_03100_));
 sky130_fd_sc_hd__a211o_1 _07890_ (.A1(_02723_),
    .A2(_03099_),
    .B1(_03100_),
    .C1(_02789_),
    .X(_03101_));
 sky130_fd_sc_hd__o2111a_1 _07891_ (.A1(_03088_),
    .A2(_03094_),
    .B1(_03096_),
    .C1(_03098_),
    .D1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__o31a_1 _07892_ (.A1(_02334_),
    .A2(_03086_),
    .A3(_03087_),
    .B1(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__o21a_1 _07893_ (.A1(_03084_),
    .A2(_03085_),
    .B1(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__inv_2 _07894_ (.A(_03104_),
    .Y(\u_decod.exe_ff_res_data_i[30] ));
 sky130_fd_sc_hd__a21o_1 _07895_ (.A1(_01079_),
    .A2(_01224_),
    .B1(_02646_),
    .X(_03105_));
 sky130_fd_sc_hd__a22o_1 _07896_ (.A1(\u_rf.reg18_q[30] ),
    .A2(_01787_),
    .B1(_02368_),
    .B2(\u_rf.reg26_q[30] ),
    .X(_03106_));
 sky130_fd_sc_hd__a221o_1 _07897_ (.A1(\u_rf.reg13_q[30] ),
    .A2(_02376_),
    .B1(_02386_),
    .B2(\u_rf.reg27_q[30] ),
    .C1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__a22o_1 _07898_ (.A1(\u_rf.reg30_q[30] ),
    .A2(_01581_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[30] ),
    .X(_03108_));
 sky130_fd_sc_hd__a221o_1 _07899_ (.A1(\u_rf.reg1_q[30] ),
    .A2(_02604_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[30] ),
    .C1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__a22o_1 _07900_ (.A1(\u_rf.reg0_q[30] ),
    .A2(_01664_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[30] ),
    .X(_03110_));
 sky130_fd_sc_hd__a221o_1 _07901_ (.A1(\u_rf.reg25_q[30] ),
    .A2(_01783_),
    .B1(_01780_),
    .B2(\u_rf.reg29_q[30] ),
    .C1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__a22o_1 _07902_ (.A1(\u_rf.reg7_q[30] ),
    .A2(_01562_),
    .B1(_02363_),
    .B2(\u_rf.reg3_q[30] ),
    .X(_03112_));
 sky130_fd_sc_hd__a221o_1 _07903_ (.A1(\u_rf.reg31_q[30] ),
    .A2(_01777_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[30] ),
    .C1(_03112_),
    .X(_03113_));
 sky130_fd_sc_hd__or4_1 _07904_ (.A(_03107_),
    .B(_03109_),
    .C(_03111_),
    .D(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__a22o_1 _07905_ (.A1(\u_rf.reg5_q[30] ),
    .A2(_02664_),
    .B1(_01610_),
    .B2(\u_rf.reg12_q[30] ),
    .X(_03115_));
 sky130_fd_sc_hd__a221o_1 _07906_ (.A1(\u_rf.reg6_q[30] ),
    .A2(_01557_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[30] ),
    .C1(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__a22o_1 _07907_ (.A1(\u_rf.reg15_q[30] ),
    .A2(_02371_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[30] ),
    .X(_03117_));
 sky130_fd_sc_hd__a221o_1 _07908_ (.A1(\u_rf.reg16_q[30] ),
    .A2(_02307_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[30] ),
    .C1(_03117_),
    .X(_03118_));
 sky130_fd_sc_hd__a22o_1 _07909_ (.A1(\u_rf.reg23_q[30] ),
    .A2(_02652_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[30] ),
    .X(_03119_));
 sky130_fd_sc_hd__a221o_1 _07910_ (.A1(\u_rf.reg9_q[30] ),
    .A2(_02360_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[30] ),
    .C1(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__a22o_1 _07911_ (.A1(\u_rf.reg24_q[30] ),
    .A2(_01784_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[30] ),
    .X(_03121_));
 sky130_fd_sc_hd__a221o_1 _07912_ (.A1(\u_rf.reg21_q[30] ),
    .A2(_02364_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[30] ),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__or4_1 _07913_ (.A(_03116_),
    .B(_03118_),
    .C(_03120_),
    .D(_03122_),
    .X(_03123_));
 sky130_fd_sc_hd__o21a_1 _07914_ (.A1(_03114_),
    .A2(_03123_),
    .B1(_02359_),
    .X(_03124_));
 sky130_fd_sc_hd__a221o_1 _07915_ (.A1(\u_decod.rf_ff_res_data_i[30] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_03105_),
    .C1(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__a21o_1 _07916_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[30] ),
    .B1(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__o31a_1 _07917_ (.A1(_03041_),
    .A2(_03042_),
    .A3(_03081_),
    .B1(_01897_),
    .X(_03127_));
 sky130_fd_sc_hd__xor2_1 _07918_ (.A(_03126_),
    .B(_03127_),
    .X(\u_decod.rs2_data_nxt[30] ));
 sky130_fd_sc_hd__a21oi_1 _07919_ (.A1(_01273_),
    .A2(_03083_),
    .B1(_01272_),
    .Y(_03128_));
 sky130_fd_sc_hd__a211o_1 _07920_ (.A1(_01273_),
    .A2(_03083_),
    .B1(_01270_),
    .C1(_01272_),
    .X(_03129_));
 sky130_fd_sc_hd__o311a_1 _07921_ (.A1(_01268_),
    .A2(_01269_),
    .A3(_03128_),
    .B1(_03129_),
    .C1(_02332_),
    .X(_03130_));
 sky130_fd_sc_hd__o21a_1 _07922_ (.A1(_01268_),
    .A2(_02244_),
    .B1(_01820_),
    .X(_03131_));
 sky130_fd_sc_hd__a2bb2o_1 _07923_ (.A1_N(_01269_),
    .A2_N(_03131_),
    .B1(_02781_),
    .B2(_01268_),
    .X(_03132_));
 sky130_fd_sc_hd__o21ai_1 _07924_ (.A1(_03130_),
    .A2(_03132_),
    .B1(_01260_),
    .Y(_03133_));
 sky130_fd_sc_hd__a21boi_1 _07925_ (.A1(_02619_),
    .A2(net57),
    .B1_N(_02618_),
    .Y(_03134_));
 sky130_fd_sc_hd__mux4_1 _07926_ (.A0(_01267_),
    .A1(_01367_),
    .A2(_01289_),
    .A3(\u_decod.rs1_data_q[7] ),
    .S0(_01469_),
    .S1(_01466_),
    .X(_03135_));
 sky130_fd_sc_hd__mux4_1 _07927_ (.A0(_02874_),
    .A1(_02964_),
    .A2(_03051_),
    .A3(_03135_),
    .S0(_01477_),
    .S1(_02685_),
    .X(_03136_));
 sky130_fd_sc_hd__nor2_1 _07928_ (.A(_02723_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__a211o_1 _07929_ (.A1(_02723_),
    .A2(_03093_),
    .B1(_03137_),
    .C1(_03088_),
    .X(_03138_));
 sky130_fd_sc_hd__or3b_1 _07930_ (.A(_02789_),
    .B(_03099_),
    .C_N(_01507_),
    .X(_03139_));
 sky130_fd_sc_hd__o211a_1 _07931_ (.A1(_02621_),
    .A2(_03134_),
    .B1(_03138_),
    .C1(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__o21ai_1 _07932_ (.A1(\u_decod.pc_q_o[31] ),
    .A2(_03087_),
    .B1(_01485_),
    .Y(_03141_));
 sky130_fd_sc_hd__a21o_1 _07933_ (.A1(\u_decod.pc_q_o[31] ),
    .A2(_03087_),
    .B1(_03141_),
    .X(_03142_));
 sky130_fd_sc_hd__nand3_1 _07934_ (.A(_03133_),
    .B(_03140_),
    .C(_03142_),
    .Y(\u_decod.exe_ff_res_data_i[31] ));
 sky130_fd_sc_hd__o21a_1 _07935_ (.A1(_01224_),
    .A2(_02644_),
    .B1(\u_decod.dec0.funct7[6] ),
    .X(_03143_));
 sky130_fd_sc_hd__a22o_1 _07936_ (.A1(\u_rf.reg30_q[31] ),
    .A2(_01581_),
    .B1(_02419_),
    .B2(\u_rf.reg28_q[31] ),
    .X(_03144_));
 sky130_fd_sc_hd__a221o_1 _07937_ (.A1(\u_rf.reg9_q[31] ),
    .A2(_02360_),
    .B1(_01668_),
    .B2(\u_rf.reg8_q[31] ),
    .C1(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__a22o_1 _07938_ (.A1(\u_rf.reg6_q[31] ),
    .A2(_01557_),
    .B1(_02375_),
    .B2(\u_rf.reg11_q[31] ),
    .X(_03146_));
 sky130_fd_sc_hd__a221o_1 _07939_ (.A1(\u_rf.reg23_q[31] ),
    .A2(_02652_),
    .B1(_01654_),
    .B2(\u_rf.reg22_q[31] ),
    .C1(_03146_),
    .X(_03147_));
 sky130_fd_sc_hd__a22o_1 _07940_ (.A1(\u_rf.reg27_q[31] ),
    .A2(_02386_),
    .B1(_01776_),
    .B2(\u_rf.reg2_q[31] ),
    .X(_03148_));
 sky130_fd_sc_hd__a221o_1 _07941_ (.A1(\u_rf.reg13_q[31] ),
    .A2(_02376_),
    .B1(_01787_),
    .B2(\u_rf.reg18_q[31] ),
    .C1(_03148_),
    .X(_03149_));
 sky130_fd_sc_hd__a22o_1 _07942_ (.A1(\u_rf.reg12_q[31] ),
    .A2(_01610_),
    .B1(_02697_),
    .B2(\u_rf.reg4_q[31] ),
    .X(_03150_));
 sky130_fd_sc_hd__a221o_1 _07943_ (.A1(\u_rf.reg31_q[31] ),
    .A2(_01777_),
    .B1(_02380_),
    .B2(\u_rf.reg10_q[31] ),
    .C1(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__or4_1 _07944_ (.A(_03145_),
    .B(_03147_),
    .C(_03149_),
    .D(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__a22o_1 _07945_ (.A1(\u_rf.reg26_q[31] ),
    .A2(_02368_),
    .B1(_02385_),
    .B2(\u_rf.reg20_q[31] ),
    .X(_03153_));
 sky130_fd_sc_hd__a221o_1 _07946_ (.A1(\u_rf.reg25_q[31] ),
    .A2(_01783_),
    .B1(_01784_),
    .B2(\u_rf.reg24_q[31] ),
    .C1(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__a22o_1 _07947_ (.A1(\u_rf.reg29_q[31] ),
    .A2(_01780_),
    .B1(_02364_),
    .B2(\u_rf.reg21_q[31] ),
    .X(_03155_));
 sky130_fd_sc_hd__a221o_1 _07948_ (.A1(\u_rf.reg1_q[31] ),
    .A2(_02604_),
    .B1(_02367_),
    .B2(\u_rf.reg14_q[31] ),
    .C1(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__a22o_1 _07949_ (.A1(\u_rf.reg7_q[31] ),
    .A2(_01562_),
    .B1(_02363_),
    .B2(\u_rf.reg3_q[31] ),
    .X(_03157_));
 sky130_fd_sc_hd__a221o_1 _07950_ (.A1(\u_rf.reg0_q[31] ),
    .A2(_01664_),
    .B1(_02371_),
    .B2(\u_rf.reg15_q[31] ),
    .C1(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__a22o_1 _07951_ (.A1(\u_rf.reg16_q[31] ),
    .A2(_02307_),
    .B1(_02379_),
    .B2(\u_rf.reg17_q[31] ),
    .X(_03159_));
 sky130_fd_sc_hd__a221o_1 _07952_ (.A1(\u_rf.reg5_q[31] ),
    .A2(_02664_),
    .B1(_02665_),
    .B2(\u_rf.reg19_q[31] ),
    .C1(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__or4_1 _07953_ (.A(_03154_),
    .B(_03156_),
    .C(_03158_),
    .D(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__o21a_1 _07954_ (.A1(_03152_),
    .A2(_03161_),
    .B1(_02359_),
    .X(_03162_));
 sky130_fd_sc_hd__a221o_1 _07955_ (.A1(\u_decod.rf_ff_res_data_i[31] ),
    .A2(_02358_),
    .B1(_02743_),
    .B2(_03143_),
    .C1(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__a21o_1 _07956_ (.A1(_02357_),
    .A2(\u_decod.exe_ff_res_data_i[31] ),
    .B1(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__o41a_1 _07957_ (.A1(_03041_),
    .A2(_03042_),
    .A3(_03081_),
    .A4(_03126_),
    .B1(_01897_),
    .X(_03165_));
 sky130_fd_sc_hd__xor2_1 _07958_ (.A(_03164_),
    .B(_03165_),
    .X(\u_decod.rs2_data_nxt[31] ));
 sky130_fd_sc_hd__xor2_1 _07959_ (.A(\u_decod.dec0.unsign_extension ),
    .B(_02229_),
    .X(_03166_));
 sky130_fd_sc_hd__mux2_1 _07960_ (.A0(_03165_),
    .A1(_03166_),
    .S(_03164_),
    .X(_03167_));
 sky130_fd_sc_hd__clkbuf_1 _07961_ (.A(_03167_),
    .X(\u_decod.rs2_data_nxt[32] ));
 sky130_fd_sc_hd__a41o_1 _07962_ (.A1(_01080_),
    .A2(_01071_),
    .A3(_01075_),
    .A4(_01094_),
    .B1(_01212_),
    .X(_03168_));
 sky130_fd_sc_hd__a21oi_1 _07963_ (.A1(\u_decod.dec0.funct3[1] ),
    .A2(\u_decod.dec0.funct3[2] ),
    .B1(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__inv_2 _07964_ (.A(\u_decod.dec0.instr_i[19] ),
    .Y(_03170_));
 sky130_fd_sc_hd__buf_2 _07965_ (.A(_03170_),
    .X(_03171_));
 sky130_fd_sc_hd__nor2_2 _07966_ (.A(\u_decod.dec0.instr_i[15] ),
    .B(\u_decod.dec0.instr_i[16] ),
    .Y(_03172_));
 sky130_fd_sc_hd__nor2_2 _07967_ (.A(\u_decod.dec0.instr_i[17] ),
    .B(\u_decod.dec0.instr_i[18] ),
    .Y(_03173_));
 sky130_fd_sc_hd__and3_4 _07968_ (.A(_03171_),
    .B(_03172_),
    .C(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__buf_6 _07969_ (.A(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__clkbuf_8 _07970_ (.A(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__inv_2 _07971_ (.A(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__o31a_4 _07972_ (.A1(_01204_),
    .A2(_01226_),
    .A3(_03169_),
    .B1(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__xor2_1 _07973_ (.A(\u_decod.dec0.instr_i[18] ),
    .B(\u_decod.exe_ff_rd_adr_q_i[3] ),
    .X(_03179_));
 sky130_fd_sc_hd__inv_2 _07974_ (.A(\u_decod.dec0.instr_i[15] ),
    .Y(_03180_));
 sky130_fd_sc_hd__inv_2 _07975_ (.A(\u_decod.dec0.instr_i[17] ),
    .Y(_03181_));
 sky130_fd_sc_hd__a22o_1 _07976_ (.A1(\u_decod.dec0.instr_i[16] ),
    .A2(_01521_),
    .B1(\u_decod.exe_ff_rd_adr_q_i[2] ),
    .B2(_03181_),
    .X(_03182_));
 sky130_fd_sc_hd__a221o_1 _07977_ (.A1(_03180_),
    .A2(\u_decod.exe_ff_rd_adr_q_i[0] ),
    .B1(\u_decod.exe_ff_rd_adr_q_i[4] ),
    .B2(_03171_),
    .C1(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__o22a_1 _07978_ (.A1(\u_decod.dec0.instr_i[16] ),
    .A2(_01521_),
    .B1(\u_decod.exe_ff_rd_adr_q_i[4] ),
    .B2(_03171_),
    .X(_03184_));
 sky130_fd_sc_hd__o221a_1 _07979_ (.A1(_03180_),
    .A2(\u_decod.exe_ff_rd_adr_q_i[0] ),
    .B1(\u_decod.exe_ff_rd_adr_q_i[2] ),
    .B2(_03181_),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__or4b_1 _07980_ (.A(_01257_),
    .B(_03179_),
    .C(_03183_),
    .D_N(_03185_),
    .X(_03186_));
 sky130_fd_sc_hd__inv_2 _07981_ (.A(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__buf_2 _07982_ (.A(\u_decod.dec0.instr_i[19] ),
    .X(_03188_));
 sky130_fd_sc_hd__a22o_1 _07983_ (.A1(_01542_),
    .A2(\u_decod.dec0.instr_i[16] ),
    .B1(_03181_),
    .B2(_01531_),
    .X(_03189_));
 sky130_fd_sc_hd__inv_2 _07984_ (.A(\u_decod.dec0.instr_i[16] ),
    .Y(_03190_));
 sky130_fd_sc_hd__inv_2 _07985_ (.A(\u_decod.dec0.instr_i[18] ),
    .Y(_03191_));
 sky130_fd_sc_hd__a22o_1 _07986_ (.A1(_01532_),
    .A2(\u_decod.dec0.instr_i[17] ),
    .B1(_03170_),
    .B2(\u_decod.rf_ff_rd_adr_q_i[4] ),
    .X(_03192_));
 sky130_fd_sc_hd__a221o_1 _07987_ (.A1(\u_decod.rf_ff_rd_adr_q_i[1] ),
    .A2(_03190_),
    .B1(_03191_),
    .B2(_01536_),
    .C1(_03192_),
    .X(_03193_));
 sky130_fd_sc_hd__xor2_1 _07988_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(\u_decod.dec0.instr_i[15] ),
    .X(_03194_));
 sky130_fd_sc_hd__a2111o_1 _07989_ (.A1(_01535_),
    .A2(\u_decod.dec0.instr_i[18] ),
    .B1(_01544_),
    .C1(_03193_),
    .D1(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__a211o_1 _07990_ (.A1(_01539_),
    .A2(_03188_),
    .B1(_03189_),
    .C1(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__nor2_2 _07991_ (.A(_03187_),
    .B(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__nor2_2 _07992_ (.A(_03181_),
    .B(_03191_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_2 _07993_ (.A(\u_decod.dec0.instr_i[15] ),
    .B(_03190_),
    .Y(_03199_));
 sky130_fd_sc_hd__and3_4 _07994_ (.A(_03188_),
    .B(_03198_),
    .C(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__nor2_2 _07995_ (.A(\u_decod.dec0.instr_i[17] ),
    .B(_03191_),
    .Y(_03201_));
 sky130_fd_sc_hd__and3_4 _07996_ (.A(_03171_),
    .B(_03201_),
    .C(_03199_),
    .X(_03202_));
 sky130_fd_sc_hd__and3_2 _07997_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03201_),
    .C(_03199_),
    .X(_03203_));
 sky130_fd_sc_hd__and2_1 _07998_ (.A(\u_decod.dec0.instr_i[15] ),
    .B(_03190_),
    .X(_03204_));
 sky130_fd_sc_hd__nor2_2 _07999_ (.A(_03181_),
    .B(\u_decod.dec0.instr_i[18] ),
    .Y(_03205_));
 sky130_fd_sc_hd__and3_2 _08000_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03204_),
    .C(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__a22o_1 _08001_ (.A1(\u_rf.reg26_q[31] ),
    .A2(_03203_),
    .B1(_03206_),
    .B2(\u_rf.reg21_q[31] ),
    .X(_03207_));
 sky130_fd_sc_hd__a221o_1 _08002_ (.A1(\u_rf.reg30_q[31] ),
    .A2(_03200_),
    .B1(_03202_),
    .B2(\u_rf.reg10_q[31] ),
    .C1(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__and2_2 _08003_ (.A(\u_decod.dec0.instr_i[15] ),
    .B(\u_decod.dec0.instr_i[16] ),
    .X(_03209_));
 sky130_fd_sc_hd__and3_4 _08004_ (.A(_03188_),
    .B(_03209_),
    .C(_03198_),
    .X(_03210_));
 sky130_fd_sc_hd__and3_4 _08005_ (.A(_03171_),
    .B(_03201_),
    .C(_03209_),
    .X(_03211_));
 sky130_fd_sc_hd__and3_2 _08006_ (.A(_03170_),
    .B(_03201_),
    .C(_03204_),
    .X(_03212_));
 sky130_fd_sc_hd__and3_2 _08007_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03172_),
    .C(_03205_),
    .X(_03213_));
 sky130_fd_sc_hd__a22o_1 _08008_ (.A1(\u_rf.reg9_q[31] ),
    .A2(_03212_),
    .B1(_03213_),
    .B2(\u_rf.reg20_q[31] ),
    .X(_03214_));
 sky130_fd_sc_hd__a221o_1 _08009_ (.A1(\u_rf.reg31_q[31] ),
    .A2(_03210_),
    .B1(_03211_),
    .B2(\u_rf.reg11_q[31] ),
    .C1(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__and3_2 _08010_ (.A(_03171_),
    .B(_03172_),
    .C(_03201_),
    .X(_03216_));
 sky130_fd_sc_hd__and3_4 _08011_ (.A(_03188_),
    .B(_03198_),
    .C(_03204_),
    .X(_03217_));
 sky130_fd_sc_hd__and3_2 _08012_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03199_),
    .C(_03205_),
    .X(_03218_));
 sky130_fd_sc_hd__and3_2 _08013_ (.A(_03170_),
    .B(_03173_),
    .C(_03209_),
    .X(_03219_));
 sky130_fd_sc_hd__a22o_1 _08014_ (.A1(\u_rf.reg22_q[31] ),
    .A2(_03218_),
    .B1(_03219_),
    .B2(\u_rf.reg3_q[31] ),
    .X(_03220_));
 sky130_fd_sc_hd__a221o_1 _08015_ (.A1(\u_rf.reg8_q[31] ),
    .A2(_03216_),
    .B1(_03217_),
    .B2(\u_rf.reg29_q[31] ),
    .C1(_03220_),
    .X(_03221_));
 sky130_fd_sc_hd__and3_2 _08016_ (.A(_03188_),
    .B(_03173_),
    .C(_03199_),
    .X(_03222_));
 sky130_fd_sc_hd__and3_2 _08017_ (.A(_03188_),
    .B(_03209_),
    .C(_03205_),
    .X(_03223_));
 sky130_fd_sc_hd__and3_4 _08018_ (.A(_03170_),
    .B(_03172_),
    .C(_03205_),
    .X(_03224_));
 sky130_fd_sc_hd__and3_4 _08019_ (.A(_03188_),
    .B(_03173_),
    .C(_03204_),
    .X(_03225_));
 sky130_fd_sc_hd__a22o_1 _08020_ (.A1(\u_rf.reg4_q[31] ),
    .A2(_03224_),
    .B1(_03225_),
    .B2(\u_rf.reg17_q[31] ),
    .X(_03226_));
 sky130_fd_sc_hd__a221o_1 _08021_ (.A1(\u_rf.reg18_q[31] ),
    .A2(_03222_),
    .B1(_03223_),
    .B2(\u_rf.reg23_q[31] ),
    .C1(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__or4_1 _08022_ (.A(_03208_),
    .B(_03215_),
    .C(_03221_),
    .D(_03227_),
    .X(_03228_));
 sky130_fd_sc_hd__and3_2 _08023_ (.A(_03171_),
    .B(_03209_),
    .C(_03205_),
    .X(_03229_));
 sky130_fd_sc_hd__and3_2 _08024_ (.A(_03188_),
    .B(_03201_),
    .C(_03204_),
    .X(_03230_));
 sky130_fd_sc_hd__and3_2 _08025_ (.A(_03170_),
    .B(_03173_),
    .C(_03204_),
    .X(_03231_));
 sky130_fd_sc_hd__and3_2 _08026_ (.A(_03170_),
    .B(_03198_),
    .C(_03199_),
    .X(_03232_));
 sky130_fd_sc_hd__a22o_1 _08027_ (.A1(\u_rf.reg1_q[31] ),
    .A2(_03231_),
    .B1(_03232_),
    .B2(\u_rf.reg14_q[31] ),
    .X(_03233_));
 sky130_fd_sc_hd__a221o_1 _08028_ (.A1(\u_rf.reg7_q[31] ),
    .A2(_03229_),
    .B1(_03230_),
    .B2(\u_rf.reg25_q[31] ),
    .C1(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__and3_4 _08029_ (.A(_03171_),
    .B(_03199_),
    .C(_03205_),
    .X(_03235_));
 sky130_fd_sc_hd__and3_4 _08030_ (.A(_03171_),
    .B(_03198_),
    .C(_03204_),
    .X(_03236_));
 sky130_fd_sc_hd__and3_4 _08031_ (.A(_03170_),
    .B(_03209_),
    .C(_03198_),
    .X(_03237_));
 sky130_fd_sc_hd__and3_2 _08032_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03172_),
    .C(_03201_),
    .X(_03238_));
 sky130_fd_sc_hd__a22o_1 _08033_ (.A1(\u_rf.reg15_q[31] ),
    .A2(_03237_),
    .B1(_03238_),
    .B2(\u_rf.reg24_q[31] ),
    .X(_03239_));
 sky130_fd_sc_hd__a221o_1 _08034_ (.A1(\u_rf.reg6_q[31] ),
    .A2(_03235_),
    .B1(_03236_),
    .B2(\u_rf.reg13_q[31] ),
    .C1(_03239_),
    .X(_03240_));
 sky130_fd_sc_hd__and3_2 _08035_ (.A(_03171_),
    .B(_03172_),
    .C(_03198_),
    .X(_03241_));
 sky130_fd_sc_hd__and3_2 _08036_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03172_),
    .C(_03198_),
    .X(_03242_));
 sky130_fd_sc_hd__and3_2 _08037_ (.A(_03170_),
    .B(_03173_),
    .C(_03199_),
    .X(_03243_));
 sky130_fd_sc_hd__a22o_1 _08038_ (.A1(\u_rf.reg28_q[31] ),
    .A2(_03242_),
    .B1(_03243_),
    .B2(\u_rf.reg2_q[31] ),
    .X(_03244_));
 sky130_fd_sc_hd__a221o_1 _08039_ (.A1(\u_rf.reg0_q[31] ),
    .A2(_03174_),
    .B1(_03241_),
    .B2(\u_rf.reg12_q[31] ),
    .C1(_03244_),
    .X(_03245_));
 sky130_fd_sc_hd__and3_4 _08040_ (.A(_03188_),
    .B(_03201_),
    .C(_03209_),
    .X(_03246_));
 sky130_fd_sc_hd__and3_2 _08041_ (.A(_03188_),
    .B(_03173_),
    .C(_03209_),
    .X(_03247_));
 sky130_fd_sc_hd__and3_2 _08042_ (.A(\u_decod.dec0.instr_i[19] ),
    .B(_03172_),
    .C(_03173_),
    .X(_03248_));
 sky130_fd_sc_hd__and3_2 _08043_ (.A(_03170_),
    .B(_03204_),
    .C(_03205_),
    .X(_03249_));
 sky130_fd_sc_hd__a22o_1 _08044_ (.A1(\u_rf.reg16_q[31] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u_rf.reg5_q[31] ),
    .X(_03250_));
 sky130_fd_sc_hd__a221o_1 _08045_ (.A1(\u_rf.reg27_q[31] ),
    .A2(_03246_),
    .B1(_03247_),
    .B2(\u_rf.reg19_q[31] ),
    .C1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__or4_1 _08046_ (.A(_03234_),
    .B(_03240_),
    .C(_03245_),
    .D(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__and2_4 _08047_ (.A(_03186_),
    .B(_03196_),
    .X(_03253_));
 sky130_fd_sc_hd__o21a_1 _08048_ (.A1(_03228_),
    .A2(_03252_),
    .B1(_03253_),
    .X(_03254_));
 sky130_fd_sc_hd__a221o_1 _08049_ (.A1(\u_decod.exe_ff_res_data_i[31] ),
    .A2(_03187_),
    .B1(_03197_),
    .B2(\u_decod.rf_ff_res_data_i[31] ),
    .C1(_03254_),
    .X(_03255_));
 sky130_fd_sc_hd__and2b_1 _08050_ (.A_N(\u_decod.dec0.instr_i[5] ),
    .B(_01224_),
    .X(_03256_));
 sky130_fd_sc_hd__buf_2 _08051_ (.A(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _08052_ (.A1(_03178_),
    .A2(_03255_),
    .B1(_03257_),
    .B2(\u_decod.pc0_q_i[31] ),
    .X(\u_decod.rs1_data[31] ));
 sky130_fd_sc_hd__and2b_1 _08053_ (.A_N(\u_decod.dec0.unsign_extension ),
    .B(\u_decod.rs1_data[31] ),
    .X(_03258_));
 sky130_fd_sc_hd__clkbuf_1 _08054_ (.A(_03258_),
    .X(\u_decod.rs1_data_nxt[32] ));
 sky130_fd_sc_hd__clkbuf_4 _08055_ (.A(_03257_),
    .X(_03259_));
 sky130_fd_sc_hd__buf_2 _08056_ (.A(_03187_),
    .X(_03260_));
 sky130_fd_sc_hd__buf_2 _08057_ (.A(_03197_),
    .X(_03261_));
 sky130_fd_sc_hd__buf_6 _08058_ (.A(_03222_),
    .X(_03262_));
 sky130_fd_sc_hd__buf_6 _08059_ (.A(_03223_),
    .X(_03263_));
 sky130_fd_sc_hd__clkbuf_8 _08060_ (.A(_03224_),
    .X(_03264_));
 sky130_fd_sc_hd__buf_6 _08061_ (.A(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__buf_6 _08062_ (.A(_03225_),
    .X(_03266_));
 sky130_fd_sc_hd__buf_6 _08063_ (.A(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__a22o_1 _08064_ (.A1(\u_rf.reg4_q[0] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[0] ),
    .X(_03268_));
 sky130_fd_sc_hd__a221o_1 _08065_ (.A1(\u_rf.reg18_q[0] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[0] ),
    .C1(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__clkbuf_8 _08066_ (.A(_03216_),
    .X(_03270_));
 sky130_fd_sc_hd__buf_6 _08067_ (.A(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__clkbuf_8 _08068_ (.A(_03217_),
    .X(_03272_));
 sky130_fd_sc_hd__clkbuf_8 _08069_ (.A(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__buf_6 _08070_ (.A(_03218_),
    .X(_03274_));
 sky130_fd_sc_hd__clkbuf_8 _08071_ (.A(_03274_),
    .X(_03275_));
 sky130_fd_sc_hd__clkbuf_8 _08072_ (.A(_03219_),
    .X(_03276_));
 sky130_fd_sc_hd__clkbuf_8 _08073_ (.A(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__a22o_1 _08074_ (.A1(\u_rf.reg22_q[0] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[0] ),
    .X(_03278_));
 sky130_fd_sc_hd__a221o_1 _08075_ (.A1(\u_rf.reg8_q[0] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[0] ),
    .C1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__buf_6 _08076_ (.A(_03200_),
    .X(_03280_));
 sky130_fd_sc_hd__clkbuf_8 _08077_ (.A(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__buf_6 _08078_ (.A(_03202_),
    .X(_03282_));
 sky130_fd_sc_hd__clkbuf_8 _08079_ (.A(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__buf_8 _08080_ (.A(_03203_),
    .X(_03284_));
 sky130_fd_sc_hd__clkbuf_8 _08081_ (.A(_03206_),
    .X(_03285_));
 sky130_fd_sc_hd__buf_6 _08082_ (.A(_03285_),
    .X(_03286_));
 sky130_fd_sc_hd__a22o_1 _08083_ (.A1(\u_rf.reg26_q[0] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[0] ),
    .X(_03287_));
 sky130_fd_sc_hd__a221o_1 _08084_ (.A1(\u_rf.reg30_q[0] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[0] ),
    .C1(_03287_),
    .X(_03288_));
 sky130_fd_sc_hd__clkbuf_8 _08085_ (.A(_03210_),
    .X(_03289_));
 sky130_fd_sc_hd__clkbuf_8 _08086_ (.A(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__buf_4 _08087_ (.A(_03211_),
    .X(_03291_));
 sky130_fd_sc_hd__clkbuf_8 _08088_ (.A(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__buf_6 _08089_ (.A(_03212_),
    .X(_03293_));
 sky130_fd_sc_hd__clkbuf_8 _08090_ (.A(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__buf_6 _08091_ (.A(_03213_),
    .X(_03295_));
 sky130_fd_sc_hd__clkbuf_8 _08092_ (.A(_03295_),
    .X(_03296_));
 sky130_fd_sc_hd__a22o_1 _08093_ (.A1(\u_rf.reg9_q[0] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[0] ),
    .X(_03297_));
 sky130_fd_sc_hd__a221o_1 _08094_ (.A1(\u_rf.reg31_q[0] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[0] ),
    .C1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__or4_1 _08095_ (.A(_03269_),
    .B(_03279_),
    .C(_03288_),
    .D(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__clkbuf_8 _08096_ (.A(_03237_),
    .X(_03300_));
 sky130_fd_sc_hd__buf_6 _08097_ (.A(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__clkbuf_8 _08098_ (.A(_03238_),
    .X(_03302_));
 sky130_fd_sc_hd__clkbuf_8 _08099_ (.A(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__buf_6 _08100_ (.A(_03235_),
    .X(_03304_));
 sky130_fd_sc_hd__buf_4 _08101_ (.A(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__clkbuf_8 _08102_ (.A(_03236_),
    .X(_03306_));
 sky130_fd_sc_hd__clkbuf_8 _08103_ (.A(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__a22o_1 _08104_ (.A1(\u_rf.reg6_q[0] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[0] ),
    .X(_03308_));
 sky130_fd_sc_hd__a221o_1 _08105_ (.A1(\u_rf.reg15_q[0] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[0] ),
    .C1(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__buf_6 _08106_ (.A(_03231_),
    .X(_03310_));
 sky130_fd_sc_hd__buf_8 _08107_ (.A(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__buf_6 _08108_ (.A(_03232_),
    .X(_03312_));
 sky130_fd_sc_hd__buf_6 _08109_ (.A(_03312_),
    .X(_03313_));
 sky130_fd_sc_hd__clkbuf_8 _08110_ (.A(_03229_),
    .X(_03314_));
 sky130_fd_sc_hd__clkbuf_8 _08111_ (.A(_03230_),
    .X(_03315_));
 sky130_fd_sc_hd__a22o_1 _08112_ (.A1(\u_rf.reg7_q[0] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[0] ),
    .X(_03316_));
 sky130_fd_sc_hd__a221o_1 _08113_ (.A1(\u_rf.reg1_q[0] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[0] ),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__clkbuf_8 _08114_ (.A(_03246_),
    .X(_03318_));
 sky130_fd_sc_hd__buf_4 _08115_ (.A(_03318_),
    .X(_03319_));
 sky130_fd_sc_hd__clkbuf_8 _08116_ (.A(_03247_),
    .X(_03320_));
 sky130_fd_sc_hd__buf_4 _08117_ (.A(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__clkbuf_8 _08118_ (.A(_03248_),
    .X(_03322_));
 sky130_fd_sc_hd__clkbuf_8 _08119_ (.A(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__clkbuf_8 _08120_ (.A(_03249_),
    .X(_03324_));
 sky130_fd_sc_hd__buf_6 _08121_ (.A(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__a22o_1 _08122_ (.A1(\u_rf.reg16_q[0] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[0] ),
    .X(_03326_));
 sky130_fd_sc_hd__a221o_1 _08123_ (.A1(\u_rf.reg27_q[0] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[0] ),
    .C1(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__buf_8 _08124_ (.A(_03241_),
    .X(_03328_));
 sky130_fd_sc_hd__buf_4 _08125_ (.A(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__buf_8 _08126_ (.A(_03242_),
    .X(_03330_));
 sky130_fd_sc_hd__clkbuf_8 _08127_ (.A(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__buf_8 _08128_ (.A(_03243_),
    .X(_03332_));
 sky130_fd_sc_hd__buf_6 _08129_ (.A(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__a22o_1 _08130_ (.A1(\u_rf.reg28_q[0] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[0] ),
    .X(_03334_));
 sky130_fd_sc_hd__a221o_1 _08131_ (.A1(\u_rf.reg0_q[0] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[0] ),
    .C1(_03334_),
    .X(_03335_));
 sky130_fd_sc_hd__or4_1 _08132_ (.A(_03309_),
    .B(_03317_),
    .C(_03327_),
    .D(_03335_),
    .X(_03336_));
 sky130_fd_sc_hd__clkbuf_8 _08133_ (.A(_03253_),
    .X(_03337_));
 sky130_fd_sc_hd__o21a_1 _08134_ (.A1(_03299_),
    .A2(_03336_),
    .B1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__a221o_1 _08135_ (.A1(\u_decod.exe_ff_res_data_i[0] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[0] ),
    .C1(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__clkbuf_4 _08136_ (.A(_03178_),
    .X(_03340_));
 sky130_fd_sc_hd__a22o_1 _08137_ (.A1(\u_decod.pc0_q_i[0] ),
    .A2(_03259_),
    .B1(_03339_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[0] ));
 sky130_fd_sc_hd__clkbuf_8 _08138_ (.A(_03280_),
    .X(_03341_));
 sky130_fd_sc_hd__clkbuf_8 _08139_ (.A(_03282_),
    .X(_03342_));
 sky130_fd_sc_hd__buf_8 _08140_ (.A(_03203_),
    .X(_03343_));
 sky130_fd_sc_hd__clkbuf_8 _08141_ (.A(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__clkbuf_8 _08142_ (.A(_03285_),
    .X(_03345_));
 sky130_fd_sc_hd__a22o_1 _08143_ (.A1(\u_rf.reg26_q[1] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[1] ),
    .X(_03346_));
 sky130_fd_sc_hd__a221o_1 _08144_ (.A1(\u_rf.reg30_q[1] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[1] ),
    .C1(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__clkbuf_8 _08145_ (.A(_03293_),
    .X(_03348_));
 sky130_fd_sc_hd__buf_6 _08146_ (.A(_03295_),
    .X(_03349_));
 sky130_fd_sc_hd__a22o_1 _08147_ (.A1(\u_rf.reg9_q[1] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[1] ),
    .X(_03350_));
 sky130_fd_sc_hd__a221o_1 _08148_ (.A1(\u_rf.reg31_q[1] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[1] ),
    .C1(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__clkbuf_8 _08149_ (.A(_03222_),
    .X(_03352_));
 sky130_fd_sc_hd__buf_6 _08150_ (.A(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__clkbuf_8 _08151_ (.A(_03223_),
    .X(_03354_));
 sky130_fd_sc_hd__buf_6 _08152_ (.A(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__buf_6 _08153_ (.A(_03264_),
    .X(_03356_));
 sky130_fd_sc_hd__buf_8 _08154_ (.A(_03266_),
    .X(_03357_));
 sky130_fd_sc_hd__a22o_1 _08155_ (.A1(\u_rf.reg4_q[1] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[1] ),
    .X(_03358_));
 sky130_fd_sc_hd__a221o_1 _08156_ (.A1(\u_rf.reg18_q[1] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[1] ),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__a22o_1 _08157_ (.A1(\u_rf.reg22_q[1] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[1] ),
    .X(_03360_));
 sky130_fd_sc_hd__a221o_1 _08158_ (.A1(\u_rf.reg8_q[1] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[1] ),
    .C1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__or3_1 _08159_ (.A(_03351_),
    .B(_03359_),
    .C(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__a22o_1 _08160_ (.A1(\u_rf.reg28_q[1] ),
    .A2(_03330_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[1] ),
    .X(_03363_));
 sky130_fd_sc_hd__a221o_1 _08161_ (.A1(\u_rf.reg0_q[1] ),
    .A2(_03175_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[1] ),
    .C1(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__buf_6 _08162_ (.A(_03318_),
    .X(_03365_));
 sky130_fd_sc_hd__buf_6 _08163_ (.A(_03247_),
    .X(_03366_));
 sky130_fd_sc_hd__a22o_1 _08164_ (.A1(\u_rf.reg16_q[1] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[1] ),
    .X(_03367_));
 sky130_fd_sc_hd__a221o_1 _08165_ (.A1(\u_rf.reg27_q[1] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[1] ),
    .C1(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__buf_6 _08166_ (.A(_03229_),
    .X(_03369_));
 sky130_fd_sc_hd__buf_6 _08167_ (.A(_03230_),
    .X(_03370_));
 sky130_fd_sc_hd__a22o_1 _08168_ (.A1(\u_rf.reg1_q[1] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[1] ),
    .X(_03371_));
 sky130_fd_sc_hd__a221o_1 _08169_ (.A1(\u_rf.reg7_q[1] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[1] ),
    .C1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__buf_6 _08170_ (.A(_03300_),
    .X(_03373_));
 sky130_fd_sc_hd__buf_6 _08171_ (.A(_03302_),
    .X(_03374_));
 sky130_fd_sc_hd__a22o_1 _08172_ (.A1(\u_rf.reg6_q[1] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[1] ),
    .X(_03375_));
 sky130_fd_sc_hd__a221o_1 _08173_ (.A1(\u_rf.reg15_q[1] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[1] ),
    .C1(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__or4_1 _08174_ (.A(_03364_),
    .B(_03368_),
    .C(_03372_),
    .D(_03376_),
    .X(_03377_));
 sky130_fd_sc_hd__clkbuf_8 _08175_ (.A(_03253_),
    .X(_03378_));
 sky130_fd_sc_hd__o31a_1 _08176_ (.A1(_03347_),
    .A2(_03362_),
    .A3(_03377_),
    .B1(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__a221o_1 _08177_ (.A1(\u_decod.exe_ff_res_data_i[1] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[1] ),
    .C1(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__a22o_1 _08178_ (.A1(\u_decod.pc0_q_i[1] ),
    .A2(_03259_),
    .B1(_03380_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[1] ));
 sky130_fd_sc_hd__clkbuf_4 _08179_ (.A(_03187_),
    .X(_03381_));
 sky130_fd_sc_hd__clkbuf_4 _08180_ (.A(_03197_),
    .X(_03382_));
 sky130_fd_sc_hd__a22o_1 _08181_ (.A1(\u_rf.reg28_q[2] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[2] ),
    .X(_03383_));
 sky130_fd_sc_hd__a221o_1 _08182_ (.A1(\u_rf.reg0_q[2] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[2] ),
    .C1(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__a22o_1 _08183_ (.A1(\u_rf.reg1_q[2] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[2] ),
    .X(_03385_));
 sky130_fd_sc_hd__a221o_1 _08184_ (.A1(\u_rf.reg7_q[2] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[2] ),
    .C1(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__clkbuf_8 _08185_ (.A(_03304_),
    .X(_03387_));
 sky130_fd_sc_hd__buf_6 _08186_ (.A(_03306_),
    .X(_03388_));
 sky130_fd_sc_hd__a22o_1 _08187_ (.A1(\u_rf.reg15_q[2] ),
    .A2(_03237_),
    .B1(_03238_),
    .B2(\u_rf.reg24_q[2] ),
    .X(_03389_));
 sky130_fd_sc_hd__a221o_1 _08188_ (.A1(\u_rf.reg6_q[2] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[2] ),
    .C1(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__a22o_1 _08189_ (.A1(\u_rf.reg16_q[2] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[2] ),
    .X(_03391_));
 sky130_fd_sc_hd__a221o_1 _08190_ (.A1(\u_rf.reg27_q[2] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[2] ),
    .C1(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__or3_1 _08191_ (.A(_03386_),
    .B(_03390_),
    .C(_03392_),
    .X(_03393_));
 sky130_fd_sc_hd__a22o_1 _08192_ (.A1(\u_rf.reg26_q[2] ),
    .A2(_03203_),
    .B1(_03206_),
    .B2(\u_rf.reg21_q[2] ),
    .X(_03394_));
 sky130_fd_sc_hd__a221o_1 _08193_ (.A1(\u_rf.reg30_q[2] ),
    .A2(_03280_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[2] ),
    .C1(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__a22o_1 _08194_ (.A1(\u_rf.reg9_q[2] ),
    .A2(_03212_),
    .B1(_03213_),
    .B2(\u_rf.reg20_q[2] ),
    .X(_03396_));
 sky130_fd_sc_hd__a221o_1 _08195_ (.A1(\u_rf.reg31_q[2] ),
    .A2(_03289_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[2] ),
    .C1(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__a22o_1 _08196_ (.A1(\u_rf.reg22_q[2] ),
    .A2(_03218_),
    .B1(_03219_),
    .B2(\u_rf.reg3_q[2] ),
    .X(_03398_));
 sky130_fd_sc_hd__a221o_1 _08197_ (.A1(\u_rf.reg8_q[2] ),
    .A2(_03216_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[2] ),
    .C1(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__a22o_1 _08198_ (.A1(\u_rf.reg4_q[2] ),
    .A2(_03224_),
    .B1(_03225_),
    .B2(\u_rf.reg17_q[2] ),
    .X(_03400_));
 sky130_fd_sc_hd__a221o_1 _08199_ (.A1(\u_rf.reg18_q[2] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[2] ),
    .C1(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__or4_1 _08200_ (.A(_03395_),
    .B(_03397_),
    .C(_03399_),
    .D(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__or3_1 _08201_ (.A(_03384_),
    .B(_03393_),
    .C(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__clkbuf_4 _08202_ (.A(_03253_),
    .X(_03404_));
 sky130_fd_sc_hd__a22o_1 _08203_ (.A1(\u_decod.rf_ff_res_data_i[2] ),
    .A2(_03382_),
    .B1(_03403_),
    .B2(_03404_),
    .X(_03405_));
 sky130_fd_sc_hd__a21o_1 _08204_ (.A1(\u_decod.exe_ff_res_data_i[2] ),
    .A2(_03381_),
    .B1(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__a22o_1 _08205_ (.A1(\u_decod.pc0_q_i[2] ),
    .A2(_03259_),
    .B1(_03406_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[2] ));
 sky130_fd_sc_hd__buf_6 _08206_ (.A(_03270_),
    .X(_03407_));
 sky130_fd_sc_hd__clkbuf_8 _08207_ (.A(_03272_),
    .X(_03408_));
 sky130_fd_sc_hd__buf_6 _08208_ (.A(_03218_),
    .X(_03409_));
 sky130_fd_sc_hd__buf_6 _08209_ (.A(_03219_),
    .X(_03410_));
 sky130_fd_sc_hd__a22o_1 _08210_ (.A1(\u_rf.reg22_q[3] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[3] ),
    .X(_03411_));
 sky130_fd_sc_hd__a221o_1 _08211_ (.A1(\u_rf.reg8_q[3] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[3] ),
    .C1(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__a22o_1 _08212_ (.A1(\u_rf.reg4_q[3] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[3] ),
    .X(_03413_));
 sky130_fd_sc_hd__a221o_1 _08213_ (.A1(\u_rf.reg18_q[3] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[3] ),
    .C1(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__a22o_1 _08214_ (.A1(\u_rf.reg9_q[3] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[3] ),
    .X(_03415_));
 sky130_fd_sc_hd__a221o_1 _08215_ (.A1(\u_rf.reg31_q[3] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[3] ),
    .C1(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__a22o_1 _08216_ (.A1(\u_rf.reg26_q[3] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[3] ),
    .X(_03417_));
 sky130_fd_sc_hd__a221o_1 _08217_ (.A1(\u_rf.reg30_q[3] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[3] ),
    .C1(_03417_),
    .X(_03418_));
 sky130_fd_sc_hd__or4_1 _08218_ (.A(_03412_),
    .B(_03414_),
    .C(_03416_),
    .D(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__clkbuf_8 _08219_ (.A(_03175_),
    .X(_03420_));
 sky130_fd_sc_hd__buf_6 _08220_ (.A(_03328_),
    .X(_03421_));
 sky130_fd_sc_hd__a22o_1 _08221_ (.A1(\u_rf.reg28_q[3] ),
    .A2(_03330_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[3] ),
    .X(_03422_));
 sky130_fd_sc_hd__a221o_1 _08222_ (.A1(\u_rf.reg0_q[3] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[3] ),
    .C1(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__a22o_1 _08223_ (.A1(\u_rf.reg16_q[3] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[3] ),
    .X(_03424_));
 sky130_fd_sc_hd__a221o_1 _08224_ (.A1(\u_rf.reg27_q[3] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[3] ),
    .C1(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__a22o_1 _08225_ (.A1(\u_rf.reg6_q[3] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[3] ),
    .X(_03426_));
 sky130_fd_sc_hd__a221o_1 _08226_ (.A1(\u_rf.reg15_q[3] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[3] ),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__buf_6 _08227_ (.A(_03314_),
    .X(_03428_));
 sky130_fd_sc_hd__buf_6 _08228_ (.A(_03315_),
    .X(_03429_));
 sky130_fd_sc_hd__a22o_1 _08229_ (.A1(\u_rf.reg1_q[3] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[3] ),
    .X(_03430_));
 sky130_fd_sc_hd__a221o_1 _08230_ (.A1(\u_rf.reg7_q[3] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[3] ),
    .C1(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__or4_1 _08231_ (.A(_03423_),
    .B(_03425_),
    .C(_03427_),
    .D(_03431_),
    .X(_03432_));
 sky130_fd_sc_hd__o21a_1 _08232_ (.A1(_03419_),
    .A2(_03432_),
    .B1(_03337_),
    .X(_03433_));
 sky130_fd_sc_hd__a221o_1 _08233_ (.A1(\u_decod.exe_ff_res_data_i[3] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[3] ),
    .C1(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__a22o_1 _08234_ (.A1(\u_decod.pc0_q_i[3] ),
    .A2(_03259_),
    .B1(_03434_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[3] ));
 sky130_fd_sc_hd__a22o_1 _08235_ (.A1(\u_rf.reg4_q[4] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[4] ),
    .X(_03435_));
 sky130_fd_sc_hd__a221o_1 _08236_ (.A1(\u_rf.reg18_q[4] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[4] ),
    .C1(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__a22o_1 _08237_ (.A1(\u_rf.reg22_q[4] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[4] ),
    .X(_03437_));
 sky130_fd_sc_hd__a221o_1 _08238_ (.A1(\u_rf.reg8_q[4] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[4] ),
    .C1(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__a22o_1 _08239_ (.A1(\u_rf.reg26_q[4] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[4] ),
    .X(_03439_));
 sky130_fd_sc_hd__a221o_1 _08240_ (.A1(\u_rf.reg30_q[4] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[4] ),
    .C1(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__a22o_1 _08241_ (.A1(\u_rf.reg9_q[4] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[4] ),
    .X(_03441_));
 sky130_fd_sc_hd__a221o_1 _08242_ (.A1(\u_rf.reg31_q[4] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[4] ),
    .C1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__or4_1 _08243_ (.A(_03436_),
    .B(_03438_),
    .C(_03440_),
    .D(_03442_),
    .X(_03443_));
 sky130_fd_sc_hd__a22o_1 _08244_ (.A1(\u_rf.reg6_q[4] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[4] ),
    .X(_03444_));
 sky130_fd_sc_hd__a221o_1 _08245_ (.A1(\u_rf.reg15_q[4] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[4] ),
    .C1(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_8 _08246_ (.A(_03310_),
    .X(_03446_));
 sky130_fd_sc_hd__buf_6 _08247_ (.A(_03312_),
    .X(_03447_));
 sky130_fd_sc_hd__a22o_1 _08248_ (.A1(\u_rf.reg1_q[4] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[4] ),
    .X(_03448_));
 sky130_fd_sc_hd__a221o_1 _08249_ (.A1(\u_rf.reg7_q[4] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[4] ),
    .C1(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__clkbuf_8 _08250_ (.A(_03322_),
    .X(_03450_));
 sky130_fd_sc_hd__a22o_1 _08251_ (.A1(\u_rf.reg16_q[4] ),
    .A2(_03450_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[4] ),
    .X(_03451_));
 sky130_fd_sc_hd__a221o_1 _08252_ (.A1(\u_rf.reg27_q[4] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[4] ),
    .C1(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__a22o_1 _08253_ (.A1(\u_rf.reg28_q[4] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[4] ),
    .X(_03453_));
 sky130_fd_sc_hd__a221o_1 _08254_ (.A1(\u_rf.reg0_q[4] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[4] ),
    .C1(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__or4_1 _08255_ (.A(_03445_),
    .B(_03449_),
    .C(_03452_),
    .D(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__o21a_1 _08256_ (.A1(_03443_),
    .A2(_03455_),
    .B1(_03337_),
    .X(_03456_));
 sky130_fd_sc_hd__a221o_1 _08257_ (.A1(\u_decod.exe_ff_res_data_i[4] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[4] ),
    .C1(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__a22o_1 _08258_ (.A1(\u_decod.pc0_q_i[4] ),
    .A2(_03259_),
    .B1(_03457_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[4] ));
 sky130_fd_sc_hd__a22o_1 _08259_ (.A1(\u_rf.reg12_q[5] ),
    .A2(_03241_),
    .B1(_03202_),
    .B2(\u_rf.reg10_q[5] ),
    .X(_03458_));
 sky130_fd_sc_hd__a221o_1 _08260_ (.A1(\u_rf.reg15_q[5] ),
    .A2(_03300_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[5] ),
    .C1(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__a22o_1 _08261_ (.A1(\u_rf.reg9_q[5] ),
    .A2(_03293_),
    .B1(_03216_),
    .B2(\u_rf.reg8_q[5] ),
    .X(_03460_));
 sky130_fd_sc_hd__a221o_1 _08262_ (.A1(\u_rf.reg6_q[5] ),
    .A2(_03387_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[5] ),
    .C1(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__a22o_1 _08263_ (.A1(\u_rf.reg27_q[5] ),
    .A2(_03246_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[5] ),
    .X(_03462_));
 sky130_fd_sc_hd__a221o_1 _08264_ (.A1(\u_rf.reg16_q[5] ),
    .A2(_03323_),
    .B1(_03280_),
    .B2(\u_rf.reg30_q[5] ),
    .C1(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__a22o_1 _08265_ (.A1(\u_rf.reg22_q[5] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[5] ),
    .X(_03464_));
 sky130_fd_sc_hd__a221o_1 _08266_ (.A1(\u_rf.reg11_q[5] ),
    .A2(_03291_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[5] ),
    .C1(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__or4_1 _08267_ (.A(_03459_),
    .B(_03461_),
    .C(_03463_),
    .D(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__a22o_1 _08268_ (.A1(\u_rf.reg28_q[5] ),
    .A2(_03330_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[5] ),
    .X(_03467_));
 sky130_fd_sc_hd__a221o_1 _08269_ (.A1(\u_rf.reg17_q[5] ),
    .A2(_03266_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[5] ),
    .C1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__a22o_1 _08270_ (.A1(\u_rf.reg31_q[5] ),
    .A2(_03210_),
    .B1(_03343_),
    .B2(\u_rf.reg26_q[5] ),
    .X(_03469_));
 sky130_fd_sc_hd__a221o_1 _08271_ (.A1(\u_rf.reg4_q[5] ),
    .A2(_03356_),
    .B1(_03311_),
    .B2(\u_rf.reg1_q[5] ),
    .C1(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__a22o_1 _08272_ (.A1(\u_rf.reg7_q[5] ),
    .A2(_03229_),
    .B1(_03230_),
    .B2(\u_rf.reg25_q[5] ),
    .X(_03471_));
 sky130_fd_sc_hd__a221o_1 _08273_ (.A1(\u_rf.reg24_q[5] ),
    .A2(_03302_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[5] ),
    .C1(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__a22o_1 _08274_ (.A1(\u_rf.reg0_q[5] ),
    .A2(_03174_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[5] ),
    .X(_03473_));
 sky130_fd_sc_hd__a221o_1 _08275_ (.A1(\u_rf.reg18_q[5] ),
    .A2(_03262_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[5] ),
    .C1(_03473_),
    .X(_03474_));
 sky130_fd_sc_hd__or4_1 _08276_ (.A(_03468_),
    .B(_03470_),
    .C(_03472_),
    .D(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__or2_1 _08277_ (.A(_03466_),
    .B(_03475_),
    .X(_03476_));
 sky130_fd_sc_hd__a22o_1 _08278_ (.A1(\u_decod.rf_ff_res_data_i[5] ),
    .A2(_03382_),
    .B1(_03476_),
    .B2(_03404_),
    .X(_03477_));
 sky130_fd_sc_hd__a21o_1 _08279_ (.A1(\u_decod.exe_ff_res_data_i[5] ),
    .A2(_03381_),
    .B1(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__a22o_1 _08280_ (.A1(\u_decod.pc0_q_i[5] ),
    .A2(_03259_),
    .B1(_03478_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[5] ));
 sky130_fd_sc_hd__a22o_1 _08281_ (.A1(\u_rf.reg28_q[6] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[6] ),
    .X(_03479_));
 sky130_fd_sc_hd__a221o_1 _08282_ (.A1(\u_rf.reg0_q[6] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[6] ),
    .C1(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__a22o_1 _08283_ (.A1(\u_rf.reg1_q[6] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[6] ),
    .X(_03481_));
 sky130_fd_sc_hd__a221o_1 _08284_ (.A1(\u_rf.reg7_q[6] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[6] ),
    .C1(_03481_),
    .X(_03482_));
 sky130_fd_sc_hd__a22o_1 _08285_ (.A1(\u_rf.reg6_q[6] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[6] ),
    .X(_03483_));
 sky130_fd_sc_hd__a221o_1 _08286_ (.A1(\u_rf.reg15_q[6] ),
    .A2(_03300_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[6] ),
    .C1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__a22o_1 _08287_ (.A1(\u_rf.reg16_q[6] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[6] ),
    .X(_03485_));
 sky130_fd_sc_hd__a221o_1 _08288_ (.A1(\u_rf.reg27_q[6] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[6] ),
    .C1(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__or3_1 _08289_ (.A(_03482_),
    .B(_03484_),
    .C(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__a22o_1 _08290_ (.A1(\u_rf.reg26_q[6] ),
    .A2(_03203_),
    .B1(_03206_),
    .B2(\u_rf.reg21_q[6] ),
    .X(_03488_));
 sky130_fd_sc_hd__a221o_1 _08291_ (.A1(\u_rf.reg30_q[6] ),
    .A2(_03200_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[6] ),
    .C1(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__a22o_1 _08292_ (.A1(\u_rf.reg9_q[6] ),
    .A2(_03212_),
    .B1(_03213_),
    .B2(\u_rf.reg20_q[6] ),
    .X(_03490_));
 sky130_fd_sc_hd__a221o_1 _08293_ (.A1(\u_rf.reg31_q[6] ),
    .A2(_03289_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[6] ),
    .C1(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__a22o_1 _08294_ (.A1(\u_rf.reg22_q[6] ),
    .A2(_03218_),
    .B1(_03219_),
    .B2(\u_rf.reg3_q[6] ),
    .X(_03492_));
 sky130_fd_sc_hd__a221o_1 _08295_ (.A1(\u_rf.reg8_q[6] ),
    .A2(_03216_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[6] ),
    .C1(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__a22o_1 _08296_ (.A1(\u_rf.reg4_q[6] ),
    .A2(_03224_),
    .B1(_03225_),
    .B2(\u_rf.reg17_q[6] ),
    .X(_03494_));
 sky130_fd_sc_hd__a221o_1 _08297_ (.A1(\u_rf.reg18_q[6] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[6] ),
    .C1(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__or4_1 _08298_ (.A(_03489_),
    .B(_03491_),
    .C(_03493_),
    .D(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__or3_1 _08299_ (.A(_03480_),
    .B(_03487_),
    .C(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__a22o_1 _08300_ (.A1(\u_decod.rf_ff_res_data_i[6] ),
    .A2(_03382_),
    .B1(_03497_),
    .B2(_03404_),
    .X(_03498_));
 sky130_fd_sc_hd__a21o_1 _08301_ (.A1(\u_decod.exe_ff_res_data_i[6] ),
    .A2(_03381_),
    .B1(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__a22o_1 _08302_ (.A1(\u_decod.pc0_q_i[6] ),
    .A2(_03259_),
    .B1(_03499_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[6] ));
 sky130_fd_sc_hd__a22o_1 _08303_ (.A1(\u_rf.reg22_q[7] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[7] ),
    .X(_03500_));
 sky130_fd_sc_hd__a221o_1 _08304_ (.A1(\u_rf.reg8_q[7] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[7] ),
    .C1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__a22o_1 _08305_ (.A1(\u_rf.reg4_q[7] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[7] ),
    .X(_03502_));
 sky130_fd_sc_hd__a221o_1 _08306_ (.A1(\u_rf.reg18_q[7] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[7] ),
    .C1(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__buf_6 _08307_ (.A(_03289_),
    .X(_03504_));
 sky130_fd_sc_hd__buf_8 _08308_ (.A(_03291_),
    .X(_03505_));
 sky130_fd_sc_hd__a22o_1 _08309_ (.A1(\u_rf.reg9_q[7] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[7] ),
    .X(_03506_));
 sky130_fd_sc_hd__a221o_1 _08310_ (.A1(\u_rf.reg31_q[7] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[7] ),
    .C1(_03506_),
    .X(_03507_));
 sky130_fd_sc_hd__a22o_1 _08311_ (.A1(\u_rf.reg26_q[7] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[7] ),
    .X(_03508_));
 sky130_fd_sc_hd__a221o_1 _08312_ (.A1(\u_rf.reg30_q[7] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[7] ),
    .C1(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__or4_1 _08313_ (.A(_03501_),
    .B(_03503_),
    .C(_03507_),
    .D(_03509_),
    .X(_03510_));
 sky130_fd_sc_hd__a22o_1 _08314_ (.A1(\u_rf.reg6_q[7] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[7] ),
    .X(_03511_));
 sky130_fd_sc_hd__a221o_1 _08315_ (.A1(\u_rf.reg15_q[7] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[7] ),
    .C1(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__a22o_1 _08316_ (.A1(\u_rf.reg1_q[7] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[7] ),
    .X(_03513_));
 sky130_fd_sc_hd__a221o_1 _08317_ (.A1(\u_rf.reg7_q[7] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[7] ),
    .C1(_03513_),
    .X(_03514_));
 sky130_fd_sc_hd__clkbuf_8 _08318_ (.A(_03324_),
    .X(_03515_));
 sky130_fd_sc_hd__a22o_1 _08319_ (.A1(\u_rf.reg16_q[7] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[7] ),
    .X(_03516_));
 sky130_fd_sc_hd__a221o_1 _08320_ (.A1(\u_rf.reg27_q[7] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[7] ),
    .C1(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__a22o_1 _08321_ (.A1(\u_rf.reg28_q[7] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[7] ),
    .X(_03518_));
 sky130_fd_sc_hd__a221o_1 _08322_ (.A1(\u_rf.reg0_q[7] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[7] ),
    .C1(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__or4_1 _08323_ (.A(_03512_),
    .B(_03514_),
    .C(_03517_),
    .D(_03519_),
    .X(_03520_));
 sky130_fd_sc_hd__o21a_1 _08324_ (.A1(_03510_),
    .A2(_03520_),
    .B1(_03337_),
    .X(_03521_));
 sky130_fd_sc_hd__a221o_1 _08325_ (.A1(\u_decod.exe_ff_res_data_i[7] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[7] ),
    .C1(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__a22o_1 _08326_ (.A1(\u_decod.pc0_q_i[7] ),
    .A2(_03259_),
    .B1(_03522_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[7] ));
 sky130_fd_sc_hd__a22o_1 _08327_ (.A1(\u_rf.reg4_q[8] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[8] ),
    .X(_03523_));
 sky130_fd_sc_hd__a221o_1 _08328_ (.A1(\u_rf.reg18_q[8] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[8] ),
    .C1(_03523_),
    .X(_03524_));
 sky130_fd_sc_hd__a22o_1 _08329_ (.A1(\u_rf.reg22_q[8] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[8] ),
    .X(_03525_));
 sky130_fd_sc_hd__a221o_1 _08330_ (.A1(\u_rf.reg8_q[8] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[8] ),
    .C1(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__a22o_1 _08331_ (.A1(\u_rf.reg26_q[8] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[8] ),
    .X(_03527_));
 sky130_fd_sc_hd__a221o_1 _08332_ (.A1(\u_rf.reg30_q[8] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[8] ),
    .C1(_03527_),
    .X(_03528_));
 sky130_fd_sc_hd__a22o_1 _08333_ (.A1(\u_rf.reg9_q[8] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[8] ),
    .X(_03529_));
 sky130_fd_sc_hd__a221o_1 _08334_ (.A1(\u_rf.reg31_q[8] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[8] ),
    .C1(_03529_),
    .X(_03530_));
 sky130_fd_sc_hd__or4_1 _08335_ (.A(_03524_),
    .B(_03526_),
    .C(_03528_),
    .D(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__a22o_1 _08336_ (.A1(\u_rf.reg28_q[8] ),
    .A2(_03330_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[8] ),
    .X(_03532_));
 sky130_fd_sc_hd__a221o_1 _08337_ (.A1(\u_rf.reg0_q[8] ),
    .A2(_03175_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[8] ),
    .C1(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__a22o_1 _08338_ (.A1(\u_rf.reg16_q[8] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[8] ),
    .X(_03534_));
 sky130_fd_sc_hd__a221o_1 _08339_ (.A1(\u_rf.reg27_q[8] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[8] ),
    .C1(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__a22o_1 _08340_ (.A1(\u_rf.reg6_q[8] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[8] ),
    .X(_03536_));
 sky130_fd_sc_hd__a221o_1 _08341_ (.A1(\u_rf.reg15_q[8] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[8] ),
    .C1(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__a22o_1 _08342_ (.A1(\u_rf.reg1_q[8] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[8] ),
    .X(_03538_));
 sky130_fd_sc_hd__a221o_1 _08343_ (.A1(\u_rf.reg7_q[8] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[8] ),
    .C1(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__or4_1 _08344_ (.A(_03533_),
    .B(_03535_),
    .C(_03537_),
    .D(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__o21a_1 _08345_ (.A1(_03531_),
    .A2(_03540_),
    .B1(_03337_),
    .X(_03541_));
 sky130_fd_sc_hd__a221o_1 _08346_ (.A1(\u_decod.exe_ff_res_data_i[8] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[8] ),
    .C1(_03541_),
    .X(_03542_));
 sky130_fd_sc_hd__a22o_1 _08347_ (.A1(\u_decod.pc0_q_i[8] ),
    .A2(_03259_),
    .B1(_03542_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[8] ));
 sky130_fd_sc_hd__a22o_1 _08348_ (.A1(\u_rf.reg4_q[9] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[9] ),
    .X(_03543_));
 sky130_fd_sc_hd__a221o_1 _08349_ (.A1(\u_rf.reg18_q[9] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[9] ),
    .C1(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__a22o_1 _08350_ (.A1(\u_rf.reg22_q[9] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[9] ),
    .X(_03545_));
 sky130_fd_sc_hd__a221o_1 _08351_ (.A1(\u_rf.reg8_q[9] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[9] ),
    .C1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__a22o_1 _08352_ (.A1(\u_rf.reg26_q[9] ),
    .A2(_03343_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[9] ),
    .X(_03547_));
 sky130_fd_sc_hd__a221o_1 _08353_ (.A1(\u_rf.reg30_q[9] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[9] ),
    .C1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__a22o_1 _08354_ (.A1(\u_rf.reg9_q[9] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[9] ),
    .X(_03549_));
 sky130_fd_sc_hd__a221o_1 _08355_ (.A1(\u_rf.reg31_q[9] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[9] ),
    .C1(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__or4_1 _08356_ (.A(_03544_),
    .B(_03546_),
    .C(_03548_),
    .D(_03550_),
    .X(_03551_));
 sky130_fd_sc_hd__a22o_1 _08357_ (.A1(\u_rf.reg1_q[9] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[9] ),
    .X(_03552_));
 sky130_fd_sc_hd__a221o_1 _08358_ (.A1(\u_rf.reg7_q[9] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[9] ),
    .C1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__a22o_1 _08359_ (.A1(\u_rf.reg15_q[9] ),
    .A2(_03300_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[9] ),
    .X(_03554_));
 sky130_fd_sc_hd__a221o_1 _08360_ (.A1(\u_rf.reg6_q[9] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[9] ),
    .C1(_03554_),
    .X(_03555_));
 sky130_fd_sc_hd__buf_8 _08361_ (.A(_03330_),
    .X(_03556_));
 sky130_fd_sc_hd__clkbuf_8 _08362_ (.A(_03332_),
    .X(_03557_));
 sky130_fd_sc_hd__a22o_1 _08363_ (.A1(\u_rf.reg28_q[9] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[9] ),
    .X(_03558_));
 sky130_fd_sc_hd__a221o_1 _08364_ (.A1(\u_rf.reg0_q[9] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[9] ),
    .C1(_03558_),
    .X(_03559_));
 sky130_fd_sc_hd__a22o_1 _08365_ (.A1(\u_rf.reg27_q[9] ),
    .A2(_03365_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[9] ),
    .X(_03560_));
 sky130_fd_sc_hd__a221o_1 _08366_ (.A1(\u_rf.reg16_q[9] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[9] ),
    .C1(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__or4_1 _08367_ (.A(_03553_),
    .B(_03555_),
    .C(_03559_),
    .D(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__o21a_1 _08368_ (.A1(_03551_),
    .A2(_03562_),
    .B1(_03337_),
    .X(_03563_));
 sky130_fd_sc_hd__a221o_1 _08369_ (.A1(\u_decod.exe_ff_res_data_i[9] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[9] ),
    .C1(_03563_),
    .X(_03564_));
 sky130_fd_sc_hd__a22o_1 _08370_ (.A1(\u_decod.pc0_q_i[9] ),
    .A2(_03259_),
    .B1(_03564_),
    .B2(_03340_),
    .X(\u_decod.rs1_data[9] ));
 sky130_fd_sc_hd__clkbuf_4 _08371_ (.A(_03257_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_1 _08372_ (.A1(\u_rf.reg4_q[10] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[10] ),
    .X(_03566_));
 sky130_fd_sc_hd__a221o_1 _08373_ (.A1(\u_rf.reg18_q[10] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[10] ),
    .C1(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__a22o_1 _08374_ (.A1(\u_rf.reg22_q[10] ),
    .A2(_03275_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[10] ),
    .X(_03568_));
 sky130_fd_sc_hd__a221o_1 _08375_ (.A1(\u_rf.reg8_q[10] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[10] ),
    .C1(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__a22o_1 _08376_ (.A1(\u_rf.reg30_q[10] ),
    .A2(_03280_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[10] ),
    .X(_03570_));
 sky130_fd_sc_hd__a221o_1 _08377_ (.A1(\u_rf.reg26_q[10] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[10] ),
    .C1(_03570_),
    .X(_03571_));
 sky130_fd_sc_hd__a22o_1 _08378_ (.A1(\u_rf.reg31_q[10] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[10] ),
    .X(_03572_));
 sky130_fd_sc_hd__a221o_1 _08379_ (.A1(\u_rf.reg9_q[10] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[10] ),
    .C1(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__or4_1 _08380_ (.A(_03567_),
    .B(_03569_),
    .C(_03571_),
    .D(_03573_),
    .X(_03574_));
 sky130_fd_sc_hd__a22o_1 _08381_ (.A1(\u_rf.reg6_q[10] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[10] ),
    .X(_03575_));
 sky130_fd_sc_hd__a221o_1 _08382_ (.A1(\u_rf.reg15_q[10] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[10] ),
    .C1(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__a22o_1 _08383_ (.A1(\u_rf.reg1_q[10] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[10] ),
    .X(_03577_));
 sky130_fd_sc_hd__a221o_1 _08384_ (.A1(\u_rf.reg7_q[10] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[10] ),
    .C1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__a22o_1 _08385_ (.A1(\u_rf.reg16_q[10] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[10] ),
    .X(_03579_));
 sky130_fd_sc_hd__a221o_1 _08386_ (.A1(\u_rf.reg27_q[10] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[10] ),
    .C1(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_1 _08387_ (.A1(\u_rf.reg28_q[10] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[10] ),
    .X(_03581_));
 sky130_fd_sc_hd__a221o_1 _08388_ (.A1(\u_rf.reg0_q[10] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[10] ),
    .C1(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__or4_1 _08389_ (.A(_03576_),
    .B(_03578_),
    .C(_03580_),
    .D(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__o21a_1 _08390_ (.A1(_03574_),
    .A2(_03583_),
    .B1(_03337_),
    .X(_03584_));
 sky130_fd_sc_hd__a221o_1 _08391_ (.A1(\u_decod.exe_ff_res_data_i[10] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[10] ),
    .C1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__clkbuf_4 _08392_ (.A(_03178_),
    .X(_03586_));
 sky130_fd_sc_hd__a22o_1 _08393_ (.A1(\u_decod.pc0_q_i[10] ),
    .A2(_03565_),
    .B1(_03585_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[10] ));
 sky130_fd_sc_hd__a22o_1 _08394_ (.A1(\u_rf.reg22_q[11] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[11] ),
    .X(_03587_));
 sky130_fd_sc_hd__a221o_1 _08395_ (.A1(\u_rf.reg8_q[11] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[11] ),
    .C1(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__a22o_1 _08396_ (.A1(\u_rf.reg4_q[11] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[11] ),
    .X(_03589_));
 sky130_fd_sc_hd__a221o_1 _08397_ (.A1(\u_rf.reg18_q[11] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[11] ),
    .C1(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_1 _08398_ (.A1(\u_rf.reg9_q[11] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[11] ),
    .X(_03591_));
 sky130_fd_sc_hd__a221o_1 _08399_ (.A1(\u_rf.reg31_q[11] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[11] ),
    .C1(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__a22o_1 _08400_ (.A1(\u_rf.reg26_q[11] ),
    .A2(_03284_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[11] ),
    .X(_03593_));
 sky130_fd_sc_hd__a221o_1 _08401_ (.A1(\u_rf.reg30_q[11] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[11] ),
    .C1(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__or4_1 _08402_ (.A(_03588_),
    .B(_03590_),
    .C(_03592_),
    .D(_03594_),
    .X(_03595_));
 sky130_fd_sc_hd__a22o_1 _08403_ (.A1(\u_rf.reg6_q[11] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[11] ),
    .X(_03596_));
 sky130_fd_sc_hd__a221o_1 _08404_ (.A1(\u_rf.reg15_q[11] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[11] ),
    .C1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_1 _08405_ (.A1(\u_rf.reg1_q[11] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[11] ),
    .X(_03598_));
 sky130_fd_sc_hd__a221o_1 _08406_ (.A1(\u_rf.reg7_q[11] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[11] ),
    .C1(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__a22o_1 _08407_ (.A1(\u_rf.reg16_q[11] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[11] ),
    .X(_03600_));
 sky130_fd_sc_hd__a221o_1 _08408_ (.A1(\u_rf.reg27_q[11] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[11] ),
    .C1(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__a22o_1 _08409_ (.A1(\u_rf.reg28_q[11] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[11] ),
    .X(_03602_));
 sky130_fd_sc_hd__a221o_1 _08410_ (.A1(\u_rf.reg0_q[11] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[11] ),
    .C1(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__or4_1 _08411_ (.A(_03597_),
    .B(_03599_),
    .C(_03601_),
    .D(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__o21a_2 _08412_ (.A1(_03595_),
    .A2(_03604_),
    .B1(_03337_),
    .X(_03605_));
 sky130_fd_sc_hd__a221o_2 _08413_ (.A1(\u_decod.exe_ff_res_data_i[11] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[11] ),
    .C1(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__a22o_1 _08414_ (.A1(\u_decod.pc0_q_i[11] ),
    .A2(_03565_),
    .B1(_03606_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[11] ));
 sky130_fd_sc_hd__a22o_1 _08415_ (.A1(\u_rf.reg22_q[12] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[12] ),
    .X(_03607_));
 sky130_fd_sc_hd__a221o_1 _08416_ (.A1(\u_rf.reg8_q[12] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[12] ),
    .C1(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__a22o_1 _08417_ (.A1(\u_rf.reg4_q[12] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[12] ),
    .X(_03609_));
 sky130_fd_sc_hd__a221o_1 _08418_ (.A1(\u_rf.reg18_q[12] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[12] ),
    .C1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__a22o_1 _08419_ (.A1(\u_rf.reg9_q[12] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[12] ),
    .X(_03611_));
 sky130_fd_sc_hd__a221o_1 _08420_ (.A1(\u_rf.reg31_q[12] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[12] ),
    .C1(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__a22o_1 _08421_ (.A1(\u_rf.reg26_q[12] ),
    .A2(_03284_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[12] ),
    .X(_03613_));
 sky130_fd_sc_hd__a221o_1 _08422_ (.A1(\u_rf.reg30_q[12] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[12] ),
    .C1(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__or4_1 _08423_ (.A(_03608_),
    .B(_03610_),
    .C(_03612_),
    .D(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__a22o_1 _08424_ (.A1(\u_rf.reg6_q[12] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[12] ),
    .X(_03616_));
 sky130_fd_sc_hd__a221o_1 _08425_ (.A1(\u_rf.reg15_q[12] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[12] ),
    .C1(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__a22o_1 _08426_ (.A1(\u_rf.reg1_q[12] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[12] ),
    .X(_03618_));
 sky130_fd_sc_hd__a221o_1 _08427_ (.A1(\u_rf.reg7_q[12] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[12] ),
    .C1(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__a22o_1 _08428_ (.A1(\u_rf.reg16_q[12] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[12] ),
    .X(_03620_));
 sky130_fd_sc_hd__a221o_1 _08429_ (.A1(\u_rf.reg27_q[12] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[12] ),
    .C1(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__a22o_1 _08430_ (.A1(\u_rf.reg28_q[12] ),
    .A2(_03331_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[12] ),
    .X(_03622_));
 sky130_fd_sc_hd__a221o_1 _08431_ (.A1(\u_rf.reg0_q[12] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[12] ),
    .C1(_03622_),
    .X(_03623_));
 sky130_fd_sc_hd__or4_1 _08432_ (.A(_03617_),
    .B(_03619_),
    .C(_03621_),
    .D(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__o21a_1 _08433_ (.A1(_03615_),
    .A2(_03624_),
    .B1(_03337_),
    .X(_03625_));
 sky130_fd_sc_hd__a221o_2 _08434_ (.A1(\u_decod.exe_ff_res_data_i[12] ),
    .A2(_03260_),
    .B1(_03261_),
    .B2(\u_decod.rf_ff_res_data_i[12] ),
    .C1(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__a22o_1 _08435_ (.A1(\u_decod.pc0_q_i[12] ),
    .A2(_03565_),
    .B1(_03626_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[12] ));
 sky130_fd_sc_hd__a22o_1 _08436_ (.A1(\u_rf.reg29_q[13] ),
    .A2(_03217_),
    .B1(_03213_),
    .B2(\u_rf.reg20_q[13] ),
    .X(_03627_));
 sky130_fd_sc_hd__a221o_1 _08437_ (.A1(\u_rf.reg18_q[13] ),
    .A2(_03352_),
    .B1(_03348_),
    .B2(\u_rf.reg9_q[13] ),
    .C1(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__a22o_1 _08438_ (.A1(\u_rf.reg27_q[13] ),
    .A2(_03246_),
    .B1(_03247_),
    .B2(\u_rf.reg19_q[13] ),
    .X(_03629_));
 sky130_fd_sc_hd__a221o_1 _08439_ (.A1(\u_rf.reg6_q[13] ),
    .A2(_03387_),
    .B1(_03270_),
    .B2(\u_rf.reg8_q[13] ),
    .C1(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__a22o_1 _08440_ (.A1(\u_rf.reg31_q[13] ),
    .A2(_03289_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[13] ),
    .X(_03631_));
 sky130_fd_sc_hd__a221o_1 _08441_ (.A1(\u_rf.reg16_q[13] ),
    .A2(_03323_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[13] ),
    .C1(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__a22o_1 _08442_ (.A1(\u_rf.reg12_q[13] ),
    .A2(_03241_),
    .B1(_03223_),
    .B2(\u_rf.reg23_q[13] ),
    .X(_03633_));
 sky130_fd_sc_hd__a221o_1 _08443_ (.A1(\u_rf.reg26_q[13] ),
    .A2(_03344_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[13] ),
    .C1(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__or4_1 _08444_ (.A(_03628_),
    .B(_03630_),
    .C(_03632_),
    .D(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__a22o_1 _08445_ (.A1(\u_rf.reg10_q[13] ),
    .A2(_03202_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[13] ),
    .X(_03636_));
 sky130_fd_sc_hd__a221o_1 _08446_ (.A1(\u_rf.reg22_q[13] ),
    .A2(_03275_),
    .B1(_03356_),
    .B2(\u_rf.reg4_q[13] ),
    .C1(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__a22o_1 _08447_ (.A1(\u_rf.reg7_q[13] ),
    .A2(_03229_),
    .B1(_03230_),
    .B2(\u_rf.reg25_q[13] ),
    .X(_03638_));
 sky130_fd_sc_hd__a221o_1 _08448_ (.A1(\u_rf.reg3_q[13] ),
    .A2(_03276_),
    .B1(_03556_),
    .B2(\u_rf.reg28_q[13] ),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a22o_1 _08449_ (.A1(\u_rf.reg24_q[13] ),
    .A2(_03238_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[13] ),
    .X(_03640_));
 sky130_fd_sc_hd__a221o_1 _08450_ (.A1(\u_rf.reg15_q[13] ),
    .A2(_03300_),
    .B1(_03311_),
    .B2(\u_rf.reg1_q[13] ),
    .C1(_03640_),
    .X(_03641_));
 sky130_fd_sc_hd__a22o_1 _08451_ (.A1(\u_rf.reg0_q[13] ),
    .A2(_03174_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[13] ),
    .X(_03642_));
 sky130_fd_sc_hd__a221o_1 _08452_ (.A1(\u_rf.reg30_q[13] ),
    .A2(_03280_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[13] ),
    .C1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__or4_1 _08453_ (.A(_03637_),
    .B(_03639_),
    .C(_03641_),
    .D(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__or2_1 _08454_ (.A(_03635_),
    .B(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__a22o_1 _08455_ (.A1(\u_decod.rf_ff_res_data_i[13] ),
    .A2(_03382_),
    .B1(_03645_),
    .B2(_03404_),
    .X(_03646_));
 sky130_fd_sc_hd__a21o_1 _08456_ (.A1(\u_decod.exe_ff_res_data_i[13] ),
    .A2(_03381_),
    .B1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__a22o_1 _08457_ (.A1(\u_decod.pc0_q_i[13] ),
    .A2(_03565_),
    .B1(_03647_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[13] ));
 sky130_fd_sc_hd__a22o_1 _08458_ (.A1(\u_rf.reg26_q[14] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[14] ),
    .X(_03648_));
 sky130_fd_sc_hd__a221o_1 _08459_ (.A1(\u_rf.reg30_q[14] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[14] ),
    .C1(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__a22o_1 _08460_ (.A1(\u_rf.reg31_q[14] ),
    .A2(_03210_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[14] ),
    .X(_03650_));
 sky130_fd_sc_hd__a221o_1 _08461_ (.A1(\u_rf.reg9_q[14] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[14] ),
    .C1(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__a22o_1 _08462_ (.A1(\u_rf.reg4_q[14] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[14] ),
    .X(_03652_));
 sky130_fd_sc_hd__a221o_1 _08463_ (.A1(\u_rf.reg18_q[14] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[14] ),
    .C1(_03652_),
    .X(_03653_));
 sky130_fd_sc_hd__a22o_1 _08464_ (.A1(\u_rf.reg22_q[14] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[14] ),
    .X(_03654_));
 sky130_fd_sc_hd__a221o_1 _08465_ (.A1(\u_rf.reg8_q[14] ),
    .A2(_03270_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[14] ),
    .C1(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__or3_1 _08466_ (.A(_03651_),
    .B(_03653_),
    .C(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__a22o_1 _08467_ (.A1(\u_rf.reg28_q[14] ),
    .A2(_03242_),
    .B1(_03243_),
    .B2(\u_rf.reg2_q[14] ),
    .X(_03657_));
 sky130_fd_sc_hd__a221o_1 _08468_ (.A1(\u_rf.reg0_q[14] ),
    .A2(_03175_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[14] ),
    .C1(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__a22o_1 _08469_ (.A1(\u_rf.reg16_q[14] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u_rf.reg5_q[14] ),
    .X(_03659_));
 sky130_fd_sc_hd__a221o_1 _08470_ (.A1(\u_rf.reg27_q[14] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[14] ),
    .C1(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__a22o_1 _08471_ (.A1(\u_rf.reg6_q[14] ),
    .A2(_03235_),
    .B1(_03236_),
    .B2(\u_rf.reg13_q[14] ),
    .X(_03661_));
 sky130_fd_sc_hd__a221o_1 _08472_ (.A1(\u_rf.reg15_q[14] ),
    .A2(_03300_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[14] ),
    .C1(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__a22o_1 _08473_ (.A1(\u_rf.reg1_q[14] ),
    .A2(_03231_),
    .B1(_03232_),
    .B2(\u_rf.reg14_q[14] ),
    .X(_03663_));
 sky130_fd_sc_hd__a221o_1 _08474_ (.A1(\u_rf.reg7_q[14] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[14] ),
    .C1(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__or4_1 _08475_ (.A(_03658_),
    .B(_03660_),
    .C(_03662_),
    .D(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__or3_2 _08476_ (.A(_03649_),
    .B(_03656_),
    .C(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__a22o_1 _08477_ (.A1(\u_decod.rf_ff_res_data_i[14] ),
    .A2(_03382_),
    .B1(_03666_),
    .B2(_03404_),
    .X(_03667_));
 sky130_fd_sc_hd__a21o_1 _08478_ (.A1(\u_decod.exe_ff_res_data_i[14] ),
    .A2(_03381_),
    .B1(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__a22o_1 _08479_ (.A1(\u_decod.pc0_q_i[14] ),
    .A2(_03565_),
    .B1(_03668_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[14] ));
 sky130_fd_sc_hd__clkbuf_4 _08480_ (.A(_03187_),
    .X(_03669_));
 sky130_fd_sc_hd__clkbuf_4 _08481_ (.A(_03197_),
    .X(_03670_));
 sky130_fd_sc_hd__a22o_1 _08482_ (.A1(\u_rf.reg22_q[15] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[15] ),
    .X(_03671_));
 sky130_fd_sc_hd__a221o_1 _08483_ (.A1(\u_rf.reg8_q[15] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[15] ),
    .C1(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__a22o_1 _08484_ (.A1(\u_rf.reg4_q[15] ),
    .A2(_03265_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[15] ),
    .X(_03673_));
 sky130_fd_sc_hd__a221o_1 _08485_ (.A1(\u_rf.reg18_q[15] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[15] ),
    .C1(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__a22o_1 _08486_ (.A1(\u_rf.reg9_q[15] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[15] ),
    .X(_03675_));
 sky130_fd_sc_hd__a221o_1 _08487_ (.A1(\u_rf.reg31_q[15] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[15] ),
    .C1(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__a22o_1 _08488_ (.A1(\u_rf.reg26_q[15] ),
    .A2(_03284_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[15] ),
    .X(_03677_));
 sky130_fd_sc_hd__a221o_1 _08489_ (.A1(\u_rf.reg30_q[15] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[15] ),
    .C1(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__or4_1 _08490_ (.A(_03672_),
    .B(_03674_),
    .C(_03676_),
    .D(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__a22o_1 _08491_ (.A1(\u_rf.reg1_q[15] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[15] ),
    .X(_03680_));
 sky130_fd_sc_hd__a221o_1 _08492_ (.A1(\u_rf.reg7_q[15] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[15] ),
    .C1(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_1 _08493_ (.A1(\u_rf.reg6_q[15] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[15] ),
    .X(_03682_));
 sky130_fd_sc_hd__a221o_1 _08494_ (.A1(\u_rf.reg15_q[15] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[15] ),
    .C1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__a22o_1 _08495_ (.A1(\u_rf.reg28_q[15] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[15] ),
    .X(_03684_));
 sky130_fd_sc_hd__a221o_1 _08496_ (.A1(\u_rf.reg0_q[15] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[15] ),
    .C1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__a22o_1 _08497_ (.A1(\u_rf.reg16_q[15] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[15] ),
    .X(_03686_));
 sky130_fd_sc_hd__a221o_1 _08498_ (.A1(\u_rf.reg27_q[15] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[15] ),
    .C1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__or4_1 _08499_ (.A(_03681_),
    .B(_03683_),
    .C(_03685_),
    .D(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__o21a_1 _08500_ (.A1(_03679_),
    .A2(_03688_),
    .B1(_03337_),
    .X(_03689_));
 sky130_fd_sc_hd__a221o_1 _08501_ (.A1(\u_decod.exe_ff_res_data_i[15] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[15] ),
    .C1(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__a22o_1 _08502_ (.A1(\u_decod.pc0_q_i[15] ),
    .A2(_03565_),
    .B1(_03690_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[15] ));
 sky130_fd_sc_hd__a22o_1 _08503_ (.A1(\u_rf.reg4_q[16] ),
    .A2(_03264_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[16] ),
    .X(_03691_));
 sky130_fd_sc_hd__a221o_1 _08504_ (.A1(\u_rf.reg18_q[16] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[16] ),
    .C1(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__a22o_1 _08505_ (.A1(\u_rf.reg22_q[16] ),
    .A2(_03409_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[16] ),
    .X(_03693_));
 sky130_fd_sc_hd__a221o_1 _08506_ (.A1(\u_rf.reg8_q[16] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[16] ),
    .C1(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__a22o_1 _08507_ (.A1(\u_rf.reg26_q[16] ),
    .A2(_03343_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[16] ),
    .X(_03695_));
 sky130_fd_sc_hd__a221o_1 _08508_ (.A1(\u_rf.reg30_q[16] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[16] ),
    .C1(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__a22o_1 _08509_ (.A1(\u_rf.reg9_q[16] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[16] ),
    .X(_03697_));
 sky130_fd_sc_hd__a221o_1 _08510_ (.A1(\u_rf.reg31_q[16] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[16] ),
    .C1(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__or4_1 _08511_ (.A(_03692_),
    .B(_03694_),
    .C(_03696_),
    .D(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__a22o_1 _08512_ (.A1(\u_rf.reg7_q[16] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[16] ),
    .X(_03700_));
 sky130_fd_sc_hd__a221o_1 _08513_ (.A1(\u_rf.reg1_q[16] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[16] ),
    .C1(_03700_),
    .X(_03701_));
 sky130_fd_sc_hd__a22o_1 _08514_ (.A1(\u_rf.reg6_q[16] ),
    .A2(_03305_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[16] ),
    .X(_03702_));
 sky130_fd_sc_hd__a221o_1 _08515_ (.A1(\u_rf.reg15_q[16] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[16] ),
    .C1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__a22o_1 _08516_ (.A1(\u_rf.reg16_q[16] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[16] ),
    .X(_03704_));
 sky130_fd_sc_hd__a221o_1 _08517_ (.A1(\u_rf.reg27_q[16] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[16] ),
    .C1(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__a22o_1 _08518_ (.A1(\u_rf.reg28_q[16] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[16] ),
    .X(_03706_));
 sky130_fd_sc_hd__a221o_1 _08519_ (.A1(\u_rf.reg0_q[16] ),
    .A2(_03420_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[16] ),
    .C1(_03706_),
    .X(_03707_));
 sky130_fd_sc_hd__or4_1 _08520_ (.A(_03701_),
    .B(_03703_),
    .C(_03705_),
    .D(_03707_),
    .X(_03708_));
 sky130_fd_sc_hd__o21a_2 _08521_ (.A1(_03699_),
    .A2(_03708_),
    .B1(_03378_),
    .X(_03709_));
 sky130_fd_sc_hd__a221o_1 _08522_ (.A1(\u_decod.exe_ff_res_data_i[16] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[16] ),
    .C1(_03709_),
    .X(_03710_));
 sky130_fd_sc_hd__a22o_1 _08523_ (.A1(\u_decod.pc0_q_i[16] ),
    .A2(_03565_),
    .B1(_03710_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[16] ));
 sky130_fd_sc_hd__a22o_1 _08524_ (.A1(\u_rf.reg26_q[17] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[17] ),
    .X(_03711_));
 sky130_fd_sc_hd__a221o_1 _08525_ (.A1(\u_rf.reg30_q[17] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[17] ),
    .C1(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__a22o_1 _08526_ (.A1(\u_rf.reg31_q[17] ),
    .A2(_03210_),
    .B1(_03211_),
    .B2(\u_rf.reg11_q[17] ),
    .X(_03713_));
 sky130_fd_sc_hd__a221o_1 _08527_ (.A1(\u_rf.reg9_q[17] ),
    .A2(_03348_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[17] ),
    .C1(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__a22o_1 _08528_ (.A1(\u_rf.reg4_q[17] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[17] ),
    .X(_03715_));
 sky130_fd_sc_hd__a221o_1 _08529_ (.A1(\u_rf.reg18_q[17] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[17] ),
    .C1(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__a22o_1 _08530_ (.A1(\u_rf.reg22_q[17] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[17] ),
    .X(_03717_));
 sky130_fd_sc_hd__a221o_1 _08531_ (.A1(\u_rf.reg8_q[17] ),
    .A2(_03270_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[17] ),
    .C1(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__or3_1 _08532_ (.A(_03714_),
    .B(_03716_),
    .C(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__a22o_1 _08533_ (.A1(\u_rf.reg1_q[17] ),
    .A2(_03231_),
    .B1(_03232_),
    .B2(\u_rf.reg14_q[17] ),
    .X(_03720_));
 sky130_fd_sc_hd__a221o_1 _08534_ (.A1(\u_rf.reg7_q[17] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[17] ),
    .C1(_03720_),
    .X(_03721_));
 sky130_fd_sc_hd__a22o_1 _08535_ (.A1(\u_rf.reg6_q[17] ),
    .A2(_03235_),
    .B1(_03236_),
    .B2(\u_rf.reg13_q[17] ),
    .X(_03722_));
 sky130_fd_sc_hd__a221o_1 _08536_ (.A1(\u_rf.reg15_q[17] ),
    .A2(_03237_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[17] ),
    .C1(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__a22o_1 _08537_ (.A1(\u_rf.reg28_q[17] ),
    .A2(_03242_),
    .B1(_03243_),
    .B2(\u_rf.reg2_q[17] ),
    .X(_03724_));
 sky130_fd_sc_hd__a221o_1 _08538_ (.A1(\u_rf.reg0_q[17] ),
    .A2(_03175_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[17] ),
    .C1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__a22o_1 _08539_ (.A1(\u_rf.reg16_q[17] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u_rf.reg5_q[17] ),
    .X(_03726_));
 sky130_fd_sc_hd__a221o_1 _08540_ (.A1(\u_rf.reg27_q[17] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[17] ),
    .C1(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__or4_1 _08541_ (.A(_03721_),
    .B(_03723_),
    .C(_03725_),
    .D(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__or3_2 _08542_ (.A(_03712_),
    .B(_03719_),
    .C(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__a22o_1 _08543_ (.A1(\u_decod.rf_ff_res_data_i[17] ),
    .A2(_03382_),
    .B1(_03729_),
    .B2(_03404_),
    .X(_03730_));
 sky130_fd_sc_hd__a21o_1 _08544_ (.A1(\u_decod.exe_ff_res_data_i[17] ),
    .A2(_03381_),
    .B1(_03730_),
    .X(_03731_));
 sky130_fd_sc_hd__a22o_1 _08545_ (.A1(\u_decod.pc0_q_i[17] ),
    .A2(_03565_),
    .B1(_03731_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[17] ));
 sky130_fd_sc_hd__a22o_1 _08546_ (.A1(\u_rf.reg6_q[18] ),
    .A2(_03304_),
    .B1(_03225_),
    .B2(\u_rf.reg17_q[18] ),
    .X(_03732_));
 sky130_fd_sc_hd__a221o_1 _08547_ (.A1(\u_rf.reg18_q[18] ),
    .A2(_03352_),
    .B1(_03275_),
    .B2(\u_rf.reg22_q[18] ),
    .C1(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__a22o_1 _08548_ (.A1(\u_rf.reg30_q[18] ),
    .A2(_03200_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[18] ),
    .X(_03734_));
 sky130_fd_sc_hd__a221o_1 _08549_ (.A1(\u_rf.reg7_q[18] ),
    .A2(_03314_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[18] ),
    .C1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__a22o_1 _08550_ (.A1(\u_rf.reg27_q[18] ),
    .A2(_03246_),
    .B1(_03289_),
    .B2(\u_rf.reg31_q[18] ),
    .X(_03736_));
 sky130_fd_sc_hd__a221o_1 _08551_ (.A1(\u_rf.reg16_q[18] ),
    .A2(_03323_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[18] ),
    .C1(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__a22o_1 _08552_ (.A1(\u_rf.reg28_q[18] ),
    .A2(_03330_),
    .B1(_03217_),
    .B2(\u_rf.reg29_q[18] ),
    .X(_03738_));
 sky130_fd_sc_hd__a221o_1 _08553_ (.A1(\u_rf.reg26_q[18] ),
    .A2(_03344_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[18] ),
    .C1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__or4_1 _08554_ (.A(_03733_),
    .B(_03735_),
    .C(_03737_),
    .D(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__a22o_1 _08555_ (.A1(\u_rf.reg4_q[18] ),
    .A2(_03224_),
    .B1(_03211_),
    .B2(\u_rf.reg11_q[18] ),
    .X(_03741_));
 sky130_fd_sc_hd__a221o_1 _08556_ (.A1(\u_rf.reg1_q[18] ),
    .A2(_03446_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[18] ),
    .C1(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__a22o_1 _08557_ (.A1(\u_rf.reg9_q[18] ),
    .A2(_03293_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[18] ),
    .X(_03743_));
 sky130_fd_sc_hd__a221o_1 _08558_ (.A1(\u_rf.reg19_q[18] ),
    .A2(_03320_),
    .B1(_03270_),
    .B2(\u_rf.reg8_q[18] ),
    .C1(_03743_),
    .X(_03744_));
 sky130_fd_sc_hd__a22o_1 _08559_ (.A1(\u_rf.reg15_q[18] ),
    .A2(_03237_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[18] ),
    .X(_03745_));
 sky130_fd_sc_hd__a221o_1 _08560_ (.A1(\u_rf.reg25_q[18] ),
    .A2(_03315_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[18] ),
    .C1(_03745_),
    .X(_03746_));
 sky130_fd_sc_hd__a22o_1 _08561_ (.A1(\u_rf.reg0_q[18] ),
    .A2(_03174_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[18] ),
    .X(_03747_));
 sky130_fd_sc_hd__a221o_1 _08562_ (.A1(\u_rf.reg23_q[18] ),
    .A2(_03354_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[18] ),
    .C1(_03747_),
    .X(_03748_));
 sky130_fd_sc_hd__or4_1 _08563_ (.A(_03742_),
    .B(_03744_),
    .C(_03746_),
    .D(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__or2_2 _08564_ (.A(_03740_),
    .B(_03749_),
    .X(_03750_));
 sky130_fd_sc_hd__a22o_1 _08565_ (.A1(\u_decod.rf_ff_res_data_i[18] ),
    .A2(_03382_),
    .B1(_03750_),
    .B2(_03404_),
    .X(_03751_));
 sky130_fd_sc_hd__a21o_1 _08566_ (.A1(\u_decod.exe_ff_res_data_i[18] ),
    .A2(_03381_),
    .B1(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__a22o_1 _08567_ (.A1(\u_decod.pc0_q_i[18] ),
    .A2(_03565_),
    .B1(_03752_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[18] ));
 sky130_fd_sc_hd__a22o_1 _08568_ (.A1(\u_rf.reg28_q[19] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[19] ),
    .X(_03753_));
 sky130_fd_sc_hd__a221o_1 _08569_ (.A1(\u_rf.reg0_q[19] ),
    .A2(_03176_),
    .B1(_03329_),
    .B2(\u_rf.reg12_q[19] ),
    .C1(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__a22o_1 _08570_ (.A1(\u_rf.reg18_q[19] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[19] ),
    .X(_03755_));
 sky130_fd_sc_hd__a221o_1 _08571_ (.A1(\u_rf.reg4_q[19] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[19] ),
    .C1(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__a22o_1 _08572_ (.A1(\u_rf.reg22_q[19] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[19] ),
    .X(_03757_));
 sky130_fd_sc_hd__a221o_1 _08573_ (.A1(\u_rf.reg8_q[19] ),
    .A2(_03270_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[19] ),
    .C1(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__a22o_1 _08574_ (.A1(\u_rf.reg9_q[19] ),
    .A2(_03293_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[19] ),
    .X(_03759_));
 sky130_fd_sc_hd__a221o_1 _08575_ (.A1(\u_rf.reg31_q[19] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[19] ),
    .C1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__a22o_1 _08576_ (.A1(\u_rf.reg26_q[19] ),
    .A2(_03343_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[19] ),
    .X(_03761_));
 sky130_fd_sc_hd__a221o_1 _08577_ (.A1(\u_rf.reg30_q[19] ),
    .A2(_03280_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[19] ),
    .C1(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__or4_1 _08578_ (.A(_03756_),
    .B(_03758_),
    .C(_03760_),
    .D(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__a22o_1 _08579_ (.A1(\u_rf.reg27_q[19] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[19] ),
    .X(_03764_));
 sky130_fd_sc_hd__a221o_1 _08580_ (.A1(\u_rf.reg16_q[19] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[19] ),
    .C1(_03764_),
    .X(_03765_));
 sky130_fd_sc_hd__a22o_1 _08581_ (.A1(\u_rf.reg7_q[19] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[19] ),
    .X(_03766_));
 sky130_fd_sc_hd__a221o_1 _08582_ (.A1(\u_rf.reg1_q[19] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[19] ),
    .C1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__a22o_1 _08583_ (.A1(\u_rf.reg6_q[19] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[19] ),
    .X(_03768_));
 sky130_fd_sc_hd__a221o_1 _08584_ (.A1(\u_rf.reg15_q[19] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[19] ),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__or3_1 _08585_ (.A(_03765_),
    .B(_03767_),
    .C(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__o31a_2 _08586_ (.A1(_03754_),
    .A2(_03763_),
    .A3(_03770_),
    .B1(_03253_),
    .X(_03771_));
 sky130_fd_sc_hd__a221o_1 _08587_ (.A1(\u_decod.exe_ff_res_data_i[19] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[19] ),
    .C1(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__a22o_1 _08588_ (.A1(\u_decod.pc0_q_i[19] ),
    .A2(_03565_),
    .B1(_03772_),
    .B2(_03586_),
    .X(\u_decod.rs1_data[19] ));
 sky130_fd_sc_hd__clkbuf_4 _08589_ (.A(_03257_),
    .X(_03773_));
 sky130_fd_sc_hd__a22o_1 _08590_ (.A1(\u_rf.reg4_q[20] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[20] ),
    .X(_03774_));
 sky130_fd_sc_hd__a221o_1 _08591_ (.A1(\u_rf.reg18_q[20] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[20] ),
    .C1(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__a22o_1 _08592_ (.A1(\u_rf.reg22_q[20] ),
    .A2(_03409_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[20] ),
    .X(_03776_));
 sky130_fd_sc_hd__a221o_1 _08593_ (.A1(\u_rf.reg8_q[20] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[20] ),
    .C1(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__a22o_1 _08594_ (.A1(\u_rf.reg26_q[20] ),
    .A2(_03343_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[20] ),
    .X(_03778_));
 sky130_fd_sc_hd__a221o_1 _08595_ (.A1(\u_rf.reg30_q[20] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[20] ),
    .C1(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__a22o_1 _08596_ (.A1(\u_rf.reg31_q[20] ),
    .A2(_03289_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[20] ),
    .X(_03780_));
 sky130_fd_sc_hd__a221o_1 _08597_ (.A1(\u_rf.reg9_q[20] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[20] ),
    .C1(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__or4_1 _08598_ (.A(_03775_),
    .B(_03777_),
    .C(_03779_),
    .D(_03781_),
    .X(_03782_));
 sky130_fd_sc_hd__a22o_1 _08599_ (.A1(\u_rf.reg6_q[20] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[20] ),
    .X(_03783_));
 sky130_fd_sc_hd__a221o_1 _08600_ (.A1(\u_rf.reg15_q[20] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[20] ),
    .C1(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__a22o_1 _08601_ (.A1(\u_rf.reg1_q[20] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[20] ),
    .X(_03785_));
 sky130_fd_sc_hd__a221o_1 _08602_ (.A1(\u_rf.reg7_q[20] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[20] ),
    .C1(_03785_),
    .X(_03786_));
 sky130_fd_sc_hd__a22o_1 _08603_ (.A1(\u_rf.reg16_q[20] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[20] ),
    .X(_03787_));
 sky130_fd_sc_hd__a221o_1 _08604_ (.A1(\u_rf.reg27_q[20] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[20] ),
    .C1(_03787_),
    .X(_03788_));
 sky130_fd_sc_hd__a22o_1 _08605_ (.A1(\u_rf.reg28_q[20] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[20] ),
    .X(_03789_));
 sky130_fd_sc_hd__a221o_1 _08606_ (.A1(\u_rf.reg0_q[20] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[20] ),
    .C1(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__or4_1 _08607_ (.A(_03784_),
    .B(_03786_),
    .C(_03788_),
    .D(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__o21a_1 _08608_ (.A1(_03782_),
    .A2(_03791_),
    .B1(_03378_),
    .X(_03792_));
 sky130_fd_sc_hd__a221o_1 _08609_ (.A1(\u_decod.exe_ff_res_data_i[20] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[20] ),
    .C1(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__clkbuf_4 _08610_ (.A(_03178_),
    .X(_03794_));
 sky130_fd_sc_hd__a22o_1 _08611_ (.A1(\u_decod.pc0_q_i[20] ),
    .A2(_03773_),
    .B1(_03793_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[20] ));
 sky130_fd_sc_hd__a22o_1 _08612_ (.A1(\u_rf.reg22_q[21] ),
    .A2(_03274_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[21] ),
    .X(_03795_));
 sky130_fd_sc_hd__a221o_1 _08613_ (.A1(\u_rf.reg8_q[21] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[21] ),
    .C1(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__a22o_1 _08614_ (.A1(\u_rf.reg4_q[21] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[21] ),
    .X(_03797_));
 sky130_fd_sc_hd__a221o_1 _08615_ (.A1(\u_rf.reg18_q[21] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[21] ),
    .C1(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__a22o_1 _08616_ (.A1(\u_rf.reg9_q[21] ),
    .A2(_03293_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[21] ),
    .X(_03799_));
 sky130_fd_sc_hd__a221o_1 _08617_ (.A1(\u_rf.reg31_q[21] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[21] ),
    .C1(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__a22o_1 _08618_ (.A1(\u_rf.reg26_q[21] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[21] ),
    .X(_03801_));
 sky130_fd_sc_hd__a221o_1 _08619_ (.A1(\u_rf.reg30_q[21] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[21] ),
    .C1(_03801_),
    .X(_03802_));
 sky130_fd_sc_hd__or4_1 _08620_ (.A(_03796_),
    .B(_03798_),
    .C(_03800_),
    .D(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__a22o_1 _08621_ (.A1(\u_rf.reg1_q[21] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[21] ),
    .X(_03804_));
 sky130_fd_sc_hd__a221o_1 _08622_ (.A1(\u_rf.reg7_q[21] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[21] ),
    .C1(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__a22o_1 _08623_ (.A1(\u_rf.reg6_q[21] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[21] ),
    .X(_03806_));
 sky130_fd_sc_hd__a221o_1 _08624_ (.A1(\u_rf.reg15_q[21] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[21] ),
    .C1(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__a22o_1 _08625_ (.A1(\u_rf.reg28_q[21] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[21] ),
    .X(_03808_));
 sky130_fd_sc_hd__a221o_1 _08626_ (.A1(\u_rf.reg0_q[21] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[21] ),
    .C1(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__a22o_1 _08627_ (.A1(\u_rf.reg16_q[21] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[21] ),
    .X(_03810_));
 sky130_fd_sc_hd__a221o_1 _08628_ (.A1(\u_rf.reg27_q[21] ),
    .A2(_03319_),
    .B1(_03321_),
    .B2(\u_rf.reg19_q[21] ),
    .C1(_03810_),
    .X(_03811_));
 sky130_fd_sc_hd__or4_1 _08629_ (.A(_03805_),
    .B(_03807_),
    .C(_03809_),
    .D(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__o21a_1 _08630_ (.A1(_03803_),
    .A2(_03812_),
    .B1(_03378_),
    .X(_03813_));
 sky130_fd_sc_hd__a221o_1 _08631_ (.A1(\u_decod.exe_ff_res_data_i[21] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[21] ),
    .C1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__a22o_1 _08632_ (.A1(\u_decod.pc0_q_i[21] ),
    .A2(_03773_),
    .B1(_03814_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[21] ));
 sky130_fd_sc_hd__a22o_1 _08633_ (.A1(\u_rf.reg19_q[22] ),
    .A2(_03247_),
    .B1(_03202_),
    .B2(\u_rf.reg10_q[22] ),
    .X(_03815_));
 sky130_fd_sc_hd__a221o_1 _08634_ (.A1(\u_rf.reg9_q[22] ),
    .A2(_03348_),
    .B1(_03300_),
    .B2(\u_rf.reg15_q[22] ),
    .C1(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__a22o_1 _08635_ (.A1(\u_rf.reg4_q[22] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[22] ),
    .X(_03817_));
 sky130_fd_sc_hd__a221o_1 _08636_ (.A1(\u_rf.reg16_q[22] ),
    .A2(_03323_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[22] ),
    .C1(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__a22o_1 _08637_ (.A1(\u_rf.reg29_q[22] ),
    .A2(_03217_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[22] ),
    .X(_03819_));
 sky130_fd_sc_hd__a221o_1 _08638_ (.A1(\u_rf.reg22_q[22] ),
    .A2(_03275_),
    .B1(_03270_),
    .B2(\u_rf.reg8_q[22] ),
    .C1(_03819_),
    .X(_03820_));
 sky130_fd_sc_hd__a22o_1 _08639_ (.A1(\u_rf.reg30_q[22] ),
    .A2(_03200_),
    .B1(_03330_),
    .B2(\u_rf.reg28_q[22] ),
    .X(_03821_));
 sky130_fd_sc_hd__a221o_1 _08640_ (.A1(\u_rf.reg7_q[22] ),
    .A2(_03369_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[22] ),
    .C1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__or4_1 _08641_ (.A(_03816_),
    .B(_03818_),
    .C(_03820_),
    .D(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__a22o_1 _08642_ (.A1(\u_rf.reg0_q[22] ),
    .A2(_03174_),
    .B1(_03238_),
    .B2(\u_rf.reg24_q[22] ),
    .X(_03824_));
 sky130_fd_sc_hd__a221o_1 _08643_ (.A1(\u_rf.reg25_q[22] ),
    .A2(_03315_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[22] ),
    .C1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__a22o_1 _08644_ (.A1(\u_rf.reg18_q[22] ),
    .A2(_03222_),
    .B1(_03223_),
    .B2(\u_rf.reg23_q[22] ),
    .X(_03826_));
 sky130_fd_sc_hd__a221o_1 _08645_ (.A1(\u_rf.reg6_q[22] ),
    .A2(_03387_),
    .B1(_03344_),
    .B2(\u_rf.reg26_q[22] ),
    .C1(_03826_),
    .X(_03827_));
 sky130_fd_sc_hd__a22o_1 _08646_ (.A1(\u_rf.reg31_q[22] ),
    .A2(_03289_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[22] ),
    .X(_03828_));
 sky130_fd_sc_hd__a221o_1 _08647_ (.A1(\u_rf.reg27_q[22] ),
    .A2(_03318_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[22] ),
    .C1(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__a22o_1 _08648_ (.A1(\u_rf.reg13_q[22] ),
    .A2(_03306_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[22] ),
    .X(_03830_));
 sky130_fd_sc_hd__a221o_1 _08649_ (.A1(\u_rf.reg1_q[22] ),
    .A2(_03311_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[22] ),
    .C1(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__or4_1 _08650_ (.A(_03825_),
    .B(_03827_),
    .C(_03829_),
    .D(_03831_),
    .X(_03832_));
 sky130_fd_sc_hd__or2_1 _08651_ (.A(_03823_),
    .B(_03832_),
    .X(_03833_));
 sky130_fd_sc_hd__a22o_1 _08652_ (.A1(\u_decod.rf_ff_res_data_i[22] ),
    .A2(_03382_),
    .B1(_03833_),
    .B2(_03404_),
    .X(_03834_));
 sky130_fd_sc_hd__a21o_1 _08653_ (.A1(\u_decod.exe_ff_res_data_i[22] ),
    .A2(_03381_),
    .B1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__a22o_1 _08654_ (.A1(\u_decod.pc0_q_i[22] ),
    .A2(_03773_),
    .B1(_03835_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[22] ));
 sky130_fd_sc_hd__a22o_1 _08655_ (.A1(\u_rf.reg22_q[23] ),
    .A2(_03274_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[23] ),
    .X(_03836_));
 sky130_fd_sc_hd__a221o_1 _08656_ (.A1(\u_rf.reg8_q[23] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[23] ),
    .C1(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__a22o_1 _08657_ (.A1(\u_rf.reg4_q[23] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[23] ),
    .X(_03838_));
 sky130_fd_sc_hd__a221o_1 _08658_ (.A1(\u_rf.reg18_q[23] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[23] ),
    .C1(_03838_),
    .X(_03839_));
 sky130_fd_sc_hd__a22o_1 _08659_ (.A1(\u_rf.reg9_q[23] ),
    .A2(_03293_),
    .B1(_03349_),
    .B2(\u_rf.reg20_q[23] ),
    .X(_03840_));
 sky130_fd_sc_hd__a221o_1 _08660_ (.A1(\u_rf.reg31_q[23] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[23] ),
    .C1(_03840_),
    .X(_03841_));
 sky130_fd_sc_hd__a22o_1 _08661_ (.A1(\u_rf.reg26_q[23] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[23] ),
    .X(_03842_));
 sky130_fd_sc_hd__a221o_1 _08662_ (.A1(\u_rf.reg30_q[23] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[23] ),
    .C1(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__or4_1 _08663_ (.A(_03837_),
    .B(_03839_),
    .C(_03841_),
    .D(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__a22o_1 _08664_ (.A1(\u_rf.reg6_q[23] ),
    .A2(_03304_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[23] ),
    .X(_03845_));
 sky130_fd_sc_hd__a221o_1 _08665_ (.A1(\u_rf.reg15_q[23] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[23] ),
    .C1(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__a22o_1 _08666_ (.A1(\u_rf.reg1_q[23] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[23] ),
    .X(_03847_));
 sky130_fd_sc_hd__a221o_1 _08667_ (.A1(\u_rf.reg7_q[23] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[23] ),
    .C1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__a22o_1 _08668_ (.A1(\u_rf.reg16_q[23] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[23] ),
    .X(_03849_));
 sky130_fd_sc_hd__a221o_1 _08669_ (.A1(\u_rf.reg27_q[23] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[23] ),
    .C1(_03849_),
    .X(_03850_));
 sky130_fd_sc_hd__a22o_1 _08670_ (.A1(\u_rf.reg0_q[23] ),
    .A2(_03175_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[23] ),
    .X(_03851_));
 sky130_fd_sc_hd__a221o_1 _08671_ (.A1(\u_rf.reg28_q[23] ),
    .A2(_03331_),
    .B1(_03333_),
    .B2(\u_rf.reg2_q[23] ),
    .C1(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__or4_1 _08672_ (.A(_03846_),
    .B(_03848_),
    .C(_03850_),
    .D(_03852_),
    .X(_03853_));
 sky130_fd_sc_hd__o21a_1 _08673_ (.A1(_03844_),
    .A2(_03853_),
    .B1(_03378_),
    .X(_03854_));
 sky130_fd_sc_hd__a221o_1 _08674_ (.A1(\u_decod.exe_ff_res_data_i[23] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[23] ),
    .C1(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__a22o_1 _08675_ (.A1(\u_decod.pc0_q_i[23] ),
    .A2(_03773_),
    .B1(_03855_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[23] ));
 sky130_fd_sc_hd__a22o_1 _08676_ (.A1(\u_rf.reg4_q[24] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[24] ),
    .X(_03856_));
 sky130_fd_sc_hd__a221o_1 _08677_ (.A1(\u_rf.reg18_q[24] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[24] ),
    .C1(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__a22o_1 _08678_ (.A1(\u_rf.reg22_q[24] ),
    .A2(_03409_),
    .B1(_03277_),
    .B2(\u_rf.reg3_q[24] ),
    .X(_03858_));
 sky130_fd_sc_hd__a221o_1 _08679_ (.A1(\u_rf.reg8_q[24] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[24] ),
    .C1(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__a22o_1 _08680_ (.A1(\u_rf.reg26_q[24] ),
    .A2(_03343_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[24] ),
    .X(_03860_));
 sky130_fd_sc_hd__a221o_1 _08681_ (.A1(\u_rf.reg30_q[24] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[24] ),
    .C1(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__a22o_1 _08682_ (.A1(\u_rf.reg9_q[24] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[24] ),
    .X(_03862_));
 sky130_fd_sc_hd__a221o_1 _08683_ (.A1(\u_rf.reg31_q[24] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[24] ),
    .C1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__or4_1 _08684_ (.A(_03857_),
    .B(_03859_),
    .C(_03861_),
    .D(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__a22o_1 _08685_ (.A1(\u_rf.reg28_q[24] ),
    .A2(_03330_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[24] ),
    .X(_03865_));
 sky130_fd_sc_hd__a221o_1 _08686_ (.A1(\u_rf.reg0_q[24] ),
    .A2(_03175_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[24] ),
    .C1(_03865_),
    .X(_03866_));
 sky130_fd_sc_hd__a22o_1 _08687_ (.A1(\u_rf.reg16_q[24] ),
    .A2(_03322_),
    .B1(_03324_),
    .B2(\u_rf.reg5_q[24] ),
    .X(_03867_));
 sky130_fd_sc_hd__a221o_1 _08688_ (.A1(\u_rf.reg27_q[24] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[24] ),
    .C1(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__a22o_1 _08689_ (.A1(\u_rf.reg6_q[24] ),
    .A2(_03387_),
    .B1(_03388_),
    .B2(\u_rf.reg13_q[24] ),
    .X(_03869_));
 sky130_fd_sc_hd__a221o_1 _08690_ (.A1(\u_rf.reg15_q[24] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[24] ),
    .C1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__a22o_1 _08691_ (.A1(\u_rf.reg1_q[24] ),
    .A2(_03311_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[24] ),
    .X(_03871_));
 sky130_fd_sc_hd__a221o_1 _08692_ (.A1(\u_rf.reg7_q[24] ),
    .A2(_03428_),
    .B1(_03429_),
    .B2(\u_rf.reg25_q[24] ),
    .C1(_03871_),
    .X(_03872_));
 sky130_fd_sc_hd__or4_1 _08693_ (.A(_03866_),
    .B(_03868_),
    .C(_03870_),
    .D(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__o21a_1 _08694_ (.A1(_03864_),
    .A2(_03873_),
    .B1(_03378_),
    .X(_03874_));
 sky130_fd_sc_hd__a221o_1 _08695_ (.A1(\u_decod.exe_ff_res_data_i[24] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[24] ),
    .C1(_03874_),
    .X(_03875_));
 sky130_fd_sc_hd__a22o_1 _08696_ (.A1(\u_decod.pc0_q_i[24] ),
    .A2(_03773_),
    .B1(_03875_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[24] ));
 sky130_fd_sc_hd__a22o_1 _08697_ (.A1(\u_rf.reg4_q[25] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[25] ),
    .X(_03876_));
 sky130_fd_sc_hd__a221o_1 _08698_ (.A1(\u_rf.reg18_q[25] ),
    .A2(_03262_),
    .B1(_03263_),
    .B2(\u_rf.reg23_q[25] ),
    .C1(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__a22o_1 _08699_ (.A1(\u_rf.reg22_q[25] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[25] ),
    .X(_03878_));
 sky130_fd_sc_hd__a221o_1 _08700_ (.A1(\u_rf.reg8_q[25] ),
    .A2(_03271_),
    .B1(_03273_),
    .B2(\u_rf.reg29_q[25] ),
    .C1(_03878_),
    .X(_03879_));
 sky130_fd_sc_hd__a22o_1 _08701_ (.A1(\u_rf.reg26_q[25] ),
    .A2(_03343_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[25] ),
    .X(_03880_));
 sky130_fd_sc_hd__a221o_1 _08702_ (.A1(\u_rf.reg30_q[25] ),
    .A2(_03280_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[25] ),
    .C1(_03880_),
    .X(_03881_));
 sky130_fd_sc_hd__a22o_1 _08703_ (.A1(\u_rf.reg9_q[25] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[25] ),
    .X(_03882_));
 sky130_fd_sc_hd__a221o_1 _08704_ (.A1(\u_rf.reg31_q[25] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[25] ),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__or4_1 _08705_ (.A(_03877_),
    .B(_03879_),
    .C(_03881_),
    .D(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__a22o_1 _08706_ (.A1(\u_rf.reg1_q[25] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[25] ),
    .X(_03885_));
 sky130_fd_sc_hd__a221o_1 _08707_ (.A1(\u_rf.reg7_q[25] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[25] ),
    .C1(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__a22o_1 _08708_ (.A1(\u_rf.reg6_q[25] ),
    .A2(_03305_),
    .B1(_03307_),
    .B2(\u_rf.reg13_q[25] ),
    .X(_03887_));
 sky130_fd_sc_hd__a221o_1 _08709_ (.A1(\u_rf.reg15_q[25] ),
    .A2(_03301_),
    .B1(_03303_),
    .B2(\u_rf.reg24_q[25] ),
    .C1(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__a22o_1 _08710_ (.A1(\u_rf.reg28_q[25] ),
    .A2(_03330_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[25] ),
    .X(_03889_));
 sky130_fd_sc_hd__a221o_1 _08711_ (.A1(\u_rf.reg0_q[25] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[25] ),
    .C1(_03889_),
    .X(_03890_));
 sky130_fd_sc_hd__a22o_1 _08712_ (.A1(\u_rf.reg27_q[25] ),
    .A2(_03365_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[25] ),
    .X(_03891_));
 sky130_fd_sc_hd__a221o_1 _08713_ (.A1(\u_rf.reg16_q[25] ),
    .A2(_03323_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[25] ),
    .C1(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__or4_1 _08714_ (.A(_03886_),
    .B(_03888_),
    .C(_03890_),
    .D(_03892_),
    .X(_03893_));
 sky130_fd_sc_hd__o21a_1 _08715_ (.A1(_03884_),
    .A2(_03893_),
    .B1(_03378_),
    .X(_03894_));
 sky130_fd_sc_hd__a221o_1 _08716_ (.A1(\u_decod.exe_ff_res_data_i[25] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[25] ),
    .C1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__a22o_1 _08717_ (.A1(\u_decod.pc0_q_i[25] ),
    .A2(_03773_),
    .B1(_03895_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[25] ));
 sky130_fd_sc_hd__a22o_1 _08718_ (.A1(\u_rf.reg18_q[26] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[26] ),
    .X(_03896_));
 sky130_fd_sc_hd__a221o_1 _08719_ (.A1(\u_rf.reg4_q[26] ),
    .A2(_03356_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[26] ),
    .C1(_03896_),
    .X(_03897_));
 sky130_fd_sc_hd__a22o_1 _08720_ (.A1(\u_rf.reg22_q[26] ),
    .A2(_03409_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[26] ),
    .X(_03898_));
 sky130_fd_sc_hd__a221o_1 _08721_ (.A1(\u_rf.reg8_q[26] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[26] ),
    .C1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__a22o_1 _08722_ (.A1(\u_rf.reg26_q[26] ),
    .A2(_03343_),
    .B1(_03285_),
    .B2(\u_rf.reg21_q[26] ),
    .X(_03900_));
 sky130_fd_sc_hd__a221o_1 _08723_ (.A1(\u_rf.reg30_q[26] ),
    .A2(_03280_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[26] ),
    .C1(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__a22o_1 _08724_ (.A1(\u_rf.reg9_q[26] ),
    .A2(_03294_),
    .B1(_03296_),
    .B2(\u_rf.reg20_q[26] ),
    .X(_03902_));
 sky130_fd_sc_hd__a221o_1 _08725_ (.A1(\u_rf.reg31_q[26] ),
    .A2(_03290_),
    .B1(_03292_),
    .B2(\u_rf.reg11_q[26] ),
    .C1(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__or4_1 _08726_ (.A(_03897_),
    .B(_03899_),
    .C(_03901_),
    .D(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__a22o_1 _08727_ (.A1(\u_rf.reg6_q[26] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[26] ),
    .X(_03905_));
 sky130_fd_sc_hd__a221o_1 _08728_ (.A1(\u_rf.reg15_q[26] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[26] ),
    .C1(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__a22o_1 _08729_ (.A1(\u_rf.reg1_q[26] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[26] ),
    .X(_03907_));
 sky130_fd_sc_hd__a221o_1 _08730_ (.A1(\u_rf.reg7_q[26] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[26] ),
    .C1(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__a22o_1 _08731_ (.A1(\u_rf.reg16_q[26] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[26] ),
    .X(_03909_));
 sky130_fd_sc_hd__a221o_1 _08732_ (.A1(\u_rf.reg27_q[26] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[26] ),
    .C1(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__a22o_1 _08733_ (.A1(\u_rf.reg28_q[26] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[26] ),
    .X(_03911_));
 sky130_fd_sc_hd__a221o_1 _08734_ (.A1(\u_rf.reg0_q[26] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[26] ),
    .C1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__or4_1 _08735_ (.A(_03906_),
    .B(_03908_),
    .C(_03910_),
    .D(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__o21a_1 _08736_ (.A1(_03904_),
    .A2(_03913_),
    .B1(_03378_),
    .X(_03914_));
 sky130_fd_sc_hd__a221o_1 _08737_ (.A1(\u_decod.exe_ff_res_data_i[26] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[26] ),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a22o_1 _08738_ (.A1(\u_decod.pc0_q_i[26] ),
    .A2(_03773_),
    .B1(_03915_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[26] ));
 sky130_fd_sc_hd__a22o_1 _08739_ (.A1(\u_rf.reg22_q[27] ),
    .A2(_03274_),
    .B1(_03410_),
    .B2(\u_rf.reg3_q[27] ),
    .X(_03916_));
 sky130_fd_sc_hd__a221o_1 _08740_ (.A1(\u_rf.reg8_q[27] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[27] ),
    .C1(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__a22o_1 _08741_ (.A1(\u_rf.reg4_q[27] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[27] ),
    .X(_03918_));
 sky130_fd_sc_hd__a221o_1 _08742_ (.A1(\u_rf.reg18_q[27] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[27] ),
    .C1(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__a22o_1 _08743_ (.A1(\u_rf.reg9_q[27] ),
    .A2(_03293_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[27] ),
    .X(_03920_));
 sky130_fd_sc_hd__a221o_1 _08744_ (.A1(\u_rf.reg31_q[27] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[27] ),
    .C1(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__a22o_1 _08745_ (.A1(\u_rf.reg26_q[27] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[27] ),
    .X(_03922_));
 sky130_fd_sc_hd__a221o_1 _08746_ (.A1(\u_rf.reg30_q[27] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[27] ),
    .C1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__or4_1 _08747_ (.A(_03917_),
    .B(_03919_),
    .C(_03921_),
    .D(_03923_),
    .X(_03924_));
 sky130_fd_sc_hd__a22o_1 _08748_ (.A1(\u_rf.reg6_q[27] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[27] ),
    .X(_03925_));
 sky130_fd_sc_hd__a221o_1 _08749_ (.A1(\u_rf.reg15_q[27] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[27] ),
    .C1(_03925_),
    .X(_03926_));
 sky130_fd_sc_hd__a22o_1 _08750_ (.A1(\u_rf.reg1_q[27] ),
    .A2(_03446_),
    .B1(_03447_),
    .B2(\u_rf.reg14_q[27] ),
    .X(_03927_));
 sky130_fd_sc_hd__a221o_1 _08751_ (.A1(\u_rf.reg7_q[27] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[27] ),
    .C1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__a22o_1 _08752_ (.A1(\u_rf.reg16_q[27] ),
    .A2(_03450_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[27] ),
    .X(_03929_));
 sky130_fd_sc_hd__a221o_1 _08753_ (.A1(\u_rf.reg27_q[27] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[27] ),
    .C1(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__a22o_1 _08754_ (.A1(\u_rf.reg28_q[27] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[27] ),
    .X(_03931_));
 sky130_fd_sc_hd__a221o_1 _08755_ (.A1(\u_rf.reg0_q[27] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[27] ),
    .C1(_03931_),
    .X(_03932_));
 sky130_fd_sc_hd__or4_1 _08756_ (.A(_03926_),
    .B(_03928_),
    .C(_03930_),
    .D(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__o21a_1 _08757_ (.A1(_03924_),
    .A2(_03933_),
    .B1(_03378_),
    .X(_03934_));
 sky130_fd_sc_hd__a221o_1 _08758_ (.A1(\u_decod.exe_ff_res_data_i[27] ),
    .A2(_03669_),
    .B1(_03670_),
    .B2(\u_decod.rf_ff_res_data_i[27] ),
    .C1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__a22o_1 _08759_ (.A1(\u_decod.pc0_q_i[27] ),
    .A2(_03773_),
    .B1(_03935_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[27] ));
 sky130_fd_sc_hd__a22o_1 _08760_ (.A1(\u_rf.reg22_q[28] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[28] ),
    .X(_03936_));
 sky130_fd_sc_hd__a221o_1 _08761_ (.A1(\u_rf.reg8_q[28] ),
    .A2(_03407_),
    .B1(_03408_),
    .B2(\u_rf.reg29_q[28] ),
    .C1(_03936_),
    .X(_03937_));
 sky130_fd_sc_hd__a22o_1 _08762_ (.A1(\u_rf.reg4_q[28] ),
    .A2(_03265_),
    .B1(_03267_),
    .B2(\u_rf.reg17_q[28] ),
    .X(_03938_));
 sky130_fd_sc_hd__a221o_1 _08763_ (.A1(\u_rf.reg18_q[28] ),
    .A2(_03353_),
    .B1(_03355_),
    .B2(\u_rf.reg23_q[28] ),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_1 _08764_ (.A1(\u_rf.reg9_q[28] ),
    .A2(_03293_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[28] ),
    .X(_03940_));
 sky130_fd_sc_hd__a221o_1 _08765_ (.A1(\u_rf.reg31_q[28] ),
    .A2(_03504_),
    .B1(_03505_),
    .B2(\u_rf.reg11_q[28] ),
    .C1(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__a22o_1 _08766_ (.A1(\u_rf.reg26_q[28] ),
    .A2(_03284_),
    .B1(_03286_),
    .B2(\u_rf.reg21_q[28] ),
    .X(_03942_));
 sky130_fd_sc_hd__a221o_1 _08767_ (.A1(\u_rf.reg30_q[28] ),
    .A2(_03281_),
    .B1(_03283_),
    .B2(\u_rf.reg10_q[28] ),
    .C1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__or4_1 _08768_ (.A(_03937_),
    .B(_03939_),
    .C(_03941_),
    .D(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__a22o_1 _08769_ (.A1(\u_rf.reg6_q[28] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[28] ),
    .X(_03945_));
 sky130_fd_sc_hd__a221o_1 _08770_ (.A1(\u_rf.reg15_q[28] ),
    .A2(_03373_),
    .B1(_03374_),
    .B2(\u_rf.reg24_q[28] ),
    .C1(_03945_),
    .X(_03946_));
 sky130_fd_sc_hd__a22o_1 _08771_ (.A1(\u_rf.reg1_q[28] ),
    .A2(_03310_),
    .B1(_03312_),
    .B2(\u_rf.reg14_q[28] ),
    .X(_03947_));
 sky130_fd_sc_hd__a221o_1 _08772_ (.A1(\u_rf.reg7_q[28] ),
    .A2(_03369_),
    .B1(_03370_),
    .B2(\u_rf.reg25_q[28] ),
    .C1(_03947_),
    .X(_03948_));
 sky130_fd_sc_hd__a22o_1 _08773_ (.A1(\u_rf.reg16_q[28] ),
    .A2(_03322_),
    .B1(_03515_),
    .B2(\u_rf.reg5_q[28] ),
    .X(_03949_));
 sky130_fd_sc_hd__a221o_1 _08774_ (.A1(\u_rf.reg27_q[28] ),
    .A2(_03365_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[28] ),
    .C1(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__a22o_1 _08775_ (.A1(\u_rf.reg28_q[28] ),
    .A2(_03556_),
    .B1(_03557_),
    .B2(\u_rf.reg2_q[28] ),
    .X(_03951_));
 sky130_fd_sc_hd__a221o_1 _08776_ (.A1(\u_rf.reg0_q[28] ),
    .A2(_03420_),
    .B1(_03421_),
    .B2(\u_rf.reg12_q[28] ),
    .C1(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__or4_1 _08777_ (.A(_03946_),
    .B(_03948_),
    .C(_03950_),
    .D(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__o21a_1 _08778_ (.A1(_03944_),
    .A2(_03953_),
    .B1(_03378_),
    .X(_03954_));
 sky130_fd_sc_hd__a221o_1 _08779_ (.A1(\u_decod.exe_ff_res_data_i[28] ),
    .A2(_03187_),
    .B1(_03382_),
    .B2(\u_decod.rf_ff_res_data_i[28] ),
    .C1(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__a22o_1 _08780_ (.A1(\u_decod.pc0_q_i[28] ),
    .A2(_03773_),
    .B1(_03955_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[28] ));
 sky130_fd_sc_hd__a22o_1 _08781_ (.A1(\u_rf.reg18_q[29] ),
    .A2(_03222_),
    .B1(_03343_),
    .B2(\u_rf.reg26_q[29] ),
    .X(_03956_));
 sky130_fd_sc_hd__a221o_1 _08782_ (.A1(\u_rf.reg23_q[29] ),
    .A2(_03354_),
    .B1(_03311_),
    .B2(\u_rf.reg1_q[29] ),
    .C1(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__a22o_1 _08783_ (.A1(\u_rf.reg21_q[29] ),
    .A2(_03206_),
    .B1(_03211_),
    .B2(\u_rf.reg11_q[29] ),
    .X(_03958_));
 sky130_fd_sc_hd__a221o_1 _08784_ (.A1(\u_rf.reg28_q[29] ),
    .A2(_03556_),
    .B1(_03356_),
    .B2(\u_rf.reg4_q[29] ),
    .C1(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__a22o_1 _08785_ (.A1(\u_rf.reg31_q[29] ),
    .A2(_03289_),
    .B1(_03332_),
    .B2(\u_rf.reg2_q[29] ),
    .X(_03960_));
 sky130_fd_sc_hd__a221o_1 _08786_ (.A1(\u_rf.reg0_q[29] ),
    .A2(_03175_),
    .B1(_03357_),
    .B2(\u_rf.reg17_q[29] ),
    .C1(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__a22o_1 _08787_ (.A1(\u_rf.reg24_q[29] ),
    .A2(_03302_),
    .B1(_03314_),
    .B2(\u_rf.reg7_q[29] ),
    .X(_03962_));
 sky130_fd_sc_hd__a221o_1 _08788_ (.A1(\u_rf.reg25_q[29] ),
    .A2(_03370_),
    .B1(_03313_),
    .B2(\u_rf.reg14_q[29] ),
    .C1(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__or4_1 _08789_ (.A(_03957_),
    .B(_03959_),
    .C(_03961_),
    .D(_03963_),
    .X(_03964_));
 sky130_fd_sc_hd__a22o_1 _08790_ (.A1(\u_rf.reg6_q[29] ),
    .A2(_03304_),
    .B1(_03306_),
    .B2(\u_rf.reg13_q[29] ),
    .X(_03965_));
 sky130_fd_sc_hd__a221o_1 _08791_ (.A1(\u_rf.reg15_q[29] ),
    .A2(_03300_),
    .B1(_03328_),
    .B2(\u_rf.reg12_q[29] ),
    .C1(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__a22o_1 _08792_ (.A1(\u_rf.reg9_q[29] ),
    .A2(_03212_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[29] ),
    .X(_03967_));
 sky130_fd_sc_hd__a221o_1 _08793_ (.A1(\u_rf.reg8_q[29] ),
    .A2(_03270_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[29] ),
    .C1(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__a22o_1 _08794_ (.A1(\u_rf.reg16_q[29] ),
    .A2(_03322_),
    .B1(_03318_),
    .B2(\u_rf.reg27_q[29] ),
    .X(_03969_));
 sky130_fd_sc_hd__a221o_1 _08795_ (.A1(\u_rf.reg30_q[29] ),
    .A2(_03280_),
    .B1(_03325_),
    .B2(\u_rf.reg5_q[29] ),
    .C1(_03969_),
    .X(_03970_));
 sky130_fd_sc_hd__a22o_1 _08796_ (.A1(\u_rf.reg3_q[29] ),
    .A2(_03276_),
    .B1(_03282_),
    .B2(\u_rf.reg10_q[29] ),
    .X(_03971_));
 sky130_fd_sc_hd__a221o_1 _08797_ (.A1(\u_rf.reg22_q[29] ),
    .A2(_03275_),
    .B1(_03366_),
    .B2(\u_rf.reg19_q[29] ),
    .C1(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__or4_1 _08798_ (.A(_03966_),
    .B(_03968_),
    .C(_03970_),
    .D(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__or2_1 _08799_ (.A(_03964_),
    .B(_03973_),
    .X(_03974_));
 sky130_fd_sc_hd__a22o_1 _08800_ (.A1(\u_decod.rf_ff_res_data_i[29] ),
    .A2(_03382_),
    .B1(_03974_),
    .B2(_03404_),
    .X(_03975_));
 sky130_fd_sc_hd__a21o_1 _08801_ (.A1(\u_decod.exe_ff_res_data_i[29] ),
    .A2(_03381_),
    .B1(_03975_),
    .X(_03976_));
 sky130_fd_sc_hd__a22o_1 _08802_ (.A1(\u_decod.pc0_q_i[29] ),
    .A2(_03773_),
    .B1(_03976_),
    .B2(_03794_),
    .X(\u_decod.rs1_data[29] ));
 sky130_fd_sc_hd__a22o_1 _08803_ (.A1(\u_rf.reg26_q[30] ),
    .A2(_03344_),
    .B1(_03345_),
    .B2(\u_rf.reg21_q[30] ),
    .X(_03977_));
 sky130_fd_sc_hd__a221o_1 _08804_ (.A1(\u_rf.reg30_q[30] ),
    .A2(_03341_),
    .B1(_03342_),
    .B2(\u_rf.reg10_q[30] ),
    .C1(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__a22o_1 _08805_ (.A1(\u_rf.reg9_q[30] ),
    .A2(_03293_),
    .B1(_03295_),
    .B2(\u_rf.reg20_q[30] ),
    .X(_03979_));
 sky130_fd_sc_hd__a221o_1 _08806_ (.A1(\u_rf.reg31_q[30] ),
    .A2(_03289_),
    .B1(_03291_),
    .B2(\u_rf.reg11_q[30] ),
    .C1(_03979_),
    .X(_03980_));
 sky130_fd_sc_hd__a22o_1 _08807_ (.A1(\u_rf.reg4_q[30] ),
    .A2(_03264_),
    .B1(_03266_),
    .B2(\u_rf.reg17_q[30] ),
    .X(_03981_));
 sky130_fd_sc_hd__a221o_1 _08808_ (.A1(\u_rf.reg18_q[30] ),
    .A2(_03352_),
    .B1(_03354_),
    .B2(\u_rf.reg23_q[30] ),
    .C1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__a22o_1 _08809_ (.A1(\u_rf.reg22_q[30] ),
    .A2(_03274_),
    .B1(_03276_),
    .B2(\u_rf.reg3_q[30] ),
    .X(_03983_));
 sky130_fd_sc_hd__a221o_1 _08810_ (.A1(\u_rf.reg8_q[30] ),
    .A2(_03270_),
    .B1(_03272_),
    .B2(\u_rf.reg29_q[30] ),
    .C1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__or3_1 _08811_ (.A(_03980_),
    .B(_03982_),
    .C(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__a22o_1 _08812_ (.A1(\u_rf.reg28_q[30] ),
    .A2(_03242_),
    .B1(_03243_),
    .B2(\u_rf.reg2_q[30] ),
    .X(_03986_));
 sky130_fd_sc_hd__a221o_1 _08813_ (.A1(\u_rf.reg0_q[30] ),
    .A2(_03175_),
    .B1(_03241_),
    .B2(\u_rf.reg12_q[30] ),
    .C1(_03986_),
    .X(_03987_));
 sky130_fd_sc_hd__a22o_1 _08814_ (.A1(\u_rf.reg16_q[30] ),
    .A2(_03248_),
    .B1(_03249_),
    .B2(\u_rf.reg5_q[30] ),
    .X(_03988_));
 sky130_fd_sc_hd__a221o_1 _08815_ (.A1(\u_rf.reg27_q[30] ),
    .A2(_03318_),
    .B1(_03320_),
    .B2(\u_rf.reg19_q[30] ),
    .C1(_03988_),
    .X(_03989_));
 sky130_fd_sc_hd__a22o_1 _08816_ (.A1(\u_rf.reg6_q[30] ),
    .A2(_03235_),
    .B1(_03236_),
    .B2(\u_rf.reg13_q[30] ),
    .X(_03990_));
 sky130_fd_sc_hd__a221o_1 _08817_ (.A1(\u_rf.reg15_q[30] ),
    .A2(_03300_),
    .B1(_03302_),
    .B2(\u_rf.reg24_q[30] ),
    .C1(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__a22o_1 _08818_ (.A1(\u_rf.reg1_q[30] ),
    .A2(_03231_),
    .B1(_03232_),
    .B2(\u_rf.reg14_q[30] ),
    .X(_03992_));
 sky130_fd_sc_hd__a221o_1 _08819_ (.A1(\u_rf.reg7_q[30] ),
    .A2(_03314_),
    .B1(_03315_),
    .B2(\u_rf.reg25_q[30] ),
    .C1(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__or4_1 _08820_ (.A(_03987_),
    .B(_03989_),
    .C(_03991_),
    .D(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__or3_1 _08821_ (.A(_03978_),
    .B(_03985_),
    .C(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__a22o_1 _08822_ (.A1(\u_decod.rf_ff_res_data_i[30] ),
    .A2(_03197_),
    .B1(_03995_),
    .B2(_03404_),
    .X(_03996_));
 sky130_fd_sc_hd__a21o_1 _08823_ (.A1(\u_decod.exe_ff_res_data_i[30] ),
    .A2(_03381_),
    .B1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__a22o_1 _08824_ (.A1(\u_decod.pc0_q_i[30] ),
    .A2(_03257_),
    .B1(_03997_),
    .B2(_03178_),
    .X(\u_decod.rs1_data[30] ));
 sky130_fd_sc_hd__clkbuf_4 _08825_ (.A(_02621_),
    .X(_03998_));
 sky130_fd_sc_hd__and2_1 _08826_ (.A(\u_decod.branch_imm_q_o[1] ),
    .B(\u_decod.rs1_data_q[1] ),
    .X(_03999_));
 sky130_fd_sc_hd__a31o_1 _08827_ (.A1(\u_decod.branch_imm_q_o[0] ),
    .A2(_01061_),
    .A3(_01060_),
    .B1(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nor2_1 _08828_ (.A(\u_decod.rs1_data_q[2] ),
    .B(\u_decod.branch_imm_q_o[2] ),
    .Y(_04001_));
 sky130_fd_sc_hd__and2_1 _08829_ (.A(\u_decod.rs1_data_q[2] ),
    .B(\u_decod.branch_imm_q_o[2] ),
    .X(_04002_));
 sky130_fd_sc_hd__nor2_1 _08830_ (.A(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_1 _08831_ (.A(_04000_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nor2_1 _08832_ (.A(_03998_),
    .B(_04004_),
    .Y(net123));
 sky130_fd_sc_hd__or2_1 _08833_ (.A(\u_decod.rs1_data_q[3] ),
    .B(\u_decod.branch_imm_q_o[3] ),
    .X(_04005_));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(\u_decod.rs1_data_q[3] ),
    .B(\u_decod.branch_imm_q_o[3] ),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_04005_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__or2_1 _08836_ (.A(\u_decod.rs1_data_q[2] ),
    .B(\u_decod.branch_imm_q_o[2] ),
    .X(_04008_));
 sky130_fd_sc_hd__a311o_1 _08837_ (.A1(\u_decod.branch_imm_q_o[0] ),
    .A2(_01061_),
    .A3(_01060_),
    .B1(_04002_),
    .C1(_03999_),
    .X(_04009_));
 sky130_fd_sc_hd__and2_1 _08838_ (.A(_04008_),
    .B(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__xor2_1 _08839_ (.A(_04007_),
    .B(_04010_),
    .X(_04011_));
 sky130_fd_sc_hd__nor2_1 _08840_ (.A(_03998_),
    .B(_04011_),
    .Y(net126));
 sky130_fd_sc_hd__or2_1 _08841_ (.A(\u_decod.rs1_data_q[4] ),
    .B(\u_decod.branch_imm_q_o[4] ),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(\u_decod.rs1_data_q[4] ),
    .B(\u_decod.branch_imm_q_o[4] ),
    .Y(_04013_));
 sky130_fd_sc_hd__and2_1 _08843_ (.A(_04012_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__and2_1 _08844_ (.A(\u_decod.rs1_data_q[3] ),
    .B(\u_decod.branch_imm_q_o[3] ),
    .X(_04015_));
 sky130_fd_sc_hd__a31o_1 _08845_ (.A1(_04008_),
    .A2(_04005_),
    .A3(_04009_),
    .B1(_04015_),
    .X(_04016_));
 sky130_fd_sc_hd__xnor2_1 _08846_ (.A(_04014_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__nor2_1 _08847_ (.A(_03998_),
    .B(_04017_),
    .Y(net127));
 sky130_fd_sc_hd__nor2_1 _08848_ (.A(\u_decod.rs1_data_q[5] ),
    .B(\u_decod.branch_imm_q_o[5] ),
    .Y(_04018_));
 sky130_fd_sc_hd__and2_1 _08849_ (.A(\u_decod.rs1_data_q[5] ),
    .B(\u_decod.branch_imm_q_o[5] ),
    .X(_04019_));
 sky130_fd_sc_hd__nor2_1 _08850_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21boi_1 _08851_ (.A1(_04014_),
    .A2(_04016_),
    .B1_N(_04013_),
    .Y(_04021_));
 sky130_fd_sc_hd__xor2_1 _08852_ (.A(_04020_),
    .B(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__nor2_1 _08853_ (.A(_03998_),
    .B(_04022_),
    .Y(net128));
 sky130_fd_sc_hd__nor2_1 _08854_ (.A(\u_decod.rs1_data_q[6] ),
    .B(\u_decod.branch_imm_q_o[6] ),
    .Y(_04023_));
 sky130_fd_sc_hd__and2_1 _08855_ (.A(\u_decod.rs1_data_q[6] ),
    .B(\u_decod.branch_imm_q_o[6] ),
    .X(_04024_));
 sky130_fd_sc_hd__nor2_1 _08856_ (.A(_04023_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__or2_1 _08857_ (.A(\u_decod.rs1_data_q[5] ),
    .B(\u_decod.branch_imm_q_o[5] ),
    .X(_04026_));
 sky130_fd_sc_hd__a31o_1 _08858_ (.A1(\u_decod.rs1_data_q[4] ),
    .A2(\u_decod.branch_imm_q_o[4] ),
    .A3(_04026_),
    .B1(_04019_),
    .X(_04027_));
 sky130_fd_sc_hd__a31o_1 _08859_ (.A1(_04014_),
    .A2(_04016_),
    .A3(_04020_),
    .B1(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__xnor2_1 _08860_ (.A(_04025_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__nor2_1 _08861_ (.A(_03998_),
    .B(_04029_),
    .Y(net129));
 sky130_fd_sc_hd__nor2_1 _08862_ (.A(\u_decod.rs1_data_q[7] ),
    .B(\u_decod.branch_imm_q_o[7] ),
    .Y(_04030_));
 sky130_fd_sc_hd__and2_1 _08863_ (.A(\u_decod.rs1_data_q[7] ),
    .B(\u_decod.branch_imm_q_o[7] ),
    .X(_04031_));
 sky130_fd_sc_hd__nor2_1 _08864_ (.A(_04030_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__a21o_1 _08865_ (.A1(_04025_),
    .A2(_04028_),
    .B1(_04024_),
    .X(_04033_));
 sky130_fd_sc_hd__xnor2_1 _08866_ (.A(_04032_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__nor2_1 _08867_ (.A(_03998_),
    .B(_04034_),
    .Y(net130));
 sky130_fd_sc_hd__nor2_1 _08868_ (.A(\u_decod.rs1_data_q[8] ),
    .B(\u_decod.branch_imm_q_o[8] ),
    .Y(_04035_));
 sky130_fd_sc_hd__and2_1 _08869_ (.A(\u_decod.rs1_data_q[8] ),
    .B(\u_decod.branch_imm_q_o[8] ),
    .X(_04036_));
 sky130_fd_sc_hd__nor2_1 _08870_ (.A(_04035_),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__or2_1 _08871_ (.A(\u_decod.rs1_data_q[7] ),
    .B(\u_decod.branch_imm_q_o[7] ),
    .X(_04038_));
 sky130_fd_sc_hd__a31o_1 _08872_ (.A1(\u_decod.rs1_data_q[6] ),
    .A2(\u_decod.branch_imm_q_o[6] ),
    .A3(_04038_),
    .B1(_04031_),
    .X(_04039_));
 sky130_fd_sc_hd__a31o_1 _08873_ (.A1(_04025_),
    .A2(_04028_),
    .A3(_04032_),
    .B1(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__xnor2_1 _08874_ (.A(_04037_),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__nor2_1 _08875_ (.A(_03998_),
    .B(_04041_),
    .Y(net131));
 sky130_fd_sc_hd__buf_2 _08876_ (.A(_02621_),
    .X(_04042_));
 sky130_fd_sc_hd__nor2_1 _08877_ (.A(\u_decod.rs1_data_q[9] ),
    .B(\u_decod.branch_imm_q_o[9] ),
    .Y(_04043_));
 sky130_fd_sc_hd__and2_1 _08878_ (.A(\u_decod.rs1_data_q[9] ),
    .B(\u_decod.branch_imm_q_o[9] ),
    .X(_04044_));
 sky130_fd_sc_hd__nor2_1 _08879_ (.A(_04043_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__a21o_1 _08880_ (.A1(_04037_),
    .A2(_04040_),
    .B1(_04036_),
    .X(_04046_));
 sky130_fd_sc_hd__xnor2_1 _08881_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__nor2_1 _08882_ (.A(_04042_),
    .B(_04047_),
    .Y(net132));
 sky130_fd_sc_hd__nor2_1 _08883_ (.A(_01302_),
    .B(\u_decod.branch_imm_q_o[10] ),
    .Y(_04048_));
 sky130_fd_sc_hd__and2_1 _08884_ (.A(_01302_),
    .B(\u_decod.branch_imm_q_o[10] ),
    .X(_04049_));
 sky130_fd_sc_hd__nor2_1 _08885_ (.A(_04048_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__or2_1 _08886_ (.A(\u_decod.rs1_data_q[9] ),
    .B(\u_decod.branch_imm_q_o[9] ),
    .X(_04051_));
 sky130_fd_sc_hd__a31o_1 _08887_ (.A1(\u_decod.rs1_data_q[8] ),
    .A2(\u_decod.branch_imm_q_o[8] ),
    .A3(_04051_),
    .B1(_04044_),
    .X(_04052_));
 sky130_fd_sc_hd__a31o_1 _08888_ (.A1(_04037_),
    .A2(_04040_),
    .A3(_04045_),
    .B1(_04052_),
    .X(_04053_));
 sky130_fd_sc_hd__xnor2_1 _08889_ (.A(_04050_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_1 _08890_ (.A(_04042_),
    .B(_04054_),
    .Y(net102));
 sky130_fd_sc_hd__nor2_1 _08891_ (.A(\u_decod.rs1_data_q[11] ),
    .B(\u_decod.branch_imm_q_o[11] ),
    .Y(_04055_));
 sky130_fd_sc_hd__and2_1 _08892_ (.A(\u_decod.rs1_data_q[11] ),
    .B(\u_decod.branch_imm_q_o[11] ),
    .X(_04056_));
 sky130_fd_sc_hd__nor2_1 _08893_ (.A(_04055_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__a21o_1 _08894_ (.A1(_04050_),
    .A2(_04053_),
    .B1(_04049_),
    .X(_04058_));
 sky130_fd_sc_hd__xnor2_1 _08895_ (.A(_04057_),
    .B(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__nor2_1 _08896_ (.A(_04042_),
    .B(_04059_),
    .Y(net103));
 sky130_fd_sc_hd__nor2_1 _08897_ (.A(_01297_),
    .B(\u_decod.branch_imm_q_o[12] ),
    .Y(_04060_));
 sky130_fd_sc_hd__and2_1 _08898_ (.A(_01297_),
    .B(\u_decod.branch_imm_q_o[12] ),
    .X(_04061_));
 sky130_fd_sc_hd__nor2_1 _08899_ (.A(_04060_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__or2_1 _08900_ (.A(\u_decod.rs1_data_q[11] ),
    .B(\u_decod.branch_imm_q_o[11] ),
    .X(_04063_));
 sky130_fd_sc_hd__a31o_1 _08901_ (.A1(_01302_),
    .A2(\u_decod.branch_imm_q_o[10] ),
    .A3(_04063_),
    .B1(_04056_),
    .X(_04064_));
 sky130_fd_sc_hd__a31o_1 _08902_ (.A1(_04050_),
    .A2(_04053_),
    .A3(_04057_),
    .B1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__xnor2_1 _08903_ (.A(_04062_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__nor2_2 _08904_ (.A(_04042_),
    .B(_04066_),
    .Y(net104));
 sky130_fd_sc_hd__nor2_1 _08905_ (.A(\u_decod.rs1_data_q[13] ),
    .B(\u_decod.branch_imm_q_o[13] ),
    .Y(_04067_));
 sky130_fd_sc_hd__and2_1 _08906_ (.A(\u_decod.rs1_data_q[13] ),
    .B(\u_decod.branch_imm_q_o[13] ),
    .X(_04068_));
 sky130_fd_sc_hd__nor2_1 _08907_ (.A(_04067_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__a21oi_1 _08908_ (.A1(_04062_),
    .A2(_04065_),
    .B1(_04061_),
    .Y(_04070_));
 sky130_fd_sc_hd__xor2_1 _08909_ (.A(_04069_),
    .B(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__nor2_1 _08910_ (.A(_04042_),
    .B(_04071_),
    .Y(net105));
 sky130_fd_sc_hd__or2_1 _08911_ (.A(_01292_),
    .B(\u_decod.branch_imm_q_o[14] ),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _08912_ (.A(_01292_),
    .B(\u_decod.branch_imm_q_o[14] ),
    .Y(_04073_));
 sky130_fd_sc_hd__and2_1 _08913_ (.A(_04072_),
    .B(_04073_),
    .X(_04074_));
 sky130_fd_sc_hd__or2_1 _08914_ (.A(\u_decod.rs1_data_q[13] ),
    .B(\u_decod.branch_imm_q_o[13] ),
    .X(_04075_));
 sky130_fd_sc_hd__a31o_1 _08915_ (.A1(_01297_),
    .A2(\u_decod.branch_imm_q_o[12] ),
    .A3(_04075_),
    .B1(_04068_),
    .X(_04076_));
 sky130_fd_sc_hd__a31o_1 _08916_ (.A1(_04062_),
    .A2(_04065_),
    .A3(_04069_),
    .B1(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__xnor2_1 _08917_ (.A(_04074_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _08918_ (.A(_04042_),
    .B(_04078_),
    .Y(net106));
 sky130_fd_sc_hd__nor2_1 _08919_ (.A(_01289_),
    .B(\u_decod.branch_imm_q_o[15] ),
    .Y(_04079_));
 sky130_fd_sc_hd__and2_1 _08920_ (.A(_01289_),
    .B(\u_decod.branch_imm_q_o[15] ),
    .X(_04080_));
 sky130_fd_sc_hd__nor2_1 _08921_ (.A(_04079_),
    .B(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__a21boi_1 _08922_ (.A1(_04074_),
    .A2(_04077_),
    .B1_N(_04073_),
    .Y(_04082_));
 sky130_fd_sc_hd__xor2_1 _08923_ (.A(_04081_),
    .B(_04082_),
    .X(_04083_));
 sky130_fd_sc_hd__nor2_1 _08924_ (.A(_04042_),
    .B(_04083_),
    .Y(net107));
 sky130_fd_sc_hd__nor2_1 _08925_ (.A(_01388_),
    .B(\u_decod.branch_imm_q_o[16] ),
    .Y(_04084_));
 sky130_fd_sc_hd__and2_1 _08926_ (.A(_01388_),
    .B(\u_decod.branch_imm_q_o[16] ),
    .X(_04085_));
 sky130_fd_sc_hd__nor2_1 _08927_ (.A(_04084_),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__or2_1 _08928_ (.A(_01289_),
    .B(\u_decod.branch_imm_q_o[15] ),
    .X(_04087_));
 sky130_fd_sc_hd__a31o_1 _08929_ (.A1(_01292_),
    .A2(\u_decod.branch_imm_q_o[14] ),
    .A3(_04087_),
    .B1(_04080_),
    .X(_04088_));
 sky130_fd_sc_hd__a31o_1 _08930_ (.A1(_04074_),
    .A2(_04077_),
    .A3(_04081_),
    .B1(_04088_),
    .X(_04089_));
 sky130_fd_sc_hd__xnor2_1 _08931_ (.A(_04086_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__nor2_1 _08932_ (.A(_04042_),
    .B(_04090_),
    .Y(net108));
 sky130_fd_sc_hd__xor2_1 _08933_ (.A(_01380_),
    .B(\u_decod.branch_imm_q_o[17] ),
    .X(_04091_));
 sky130_fd_sc_hd__a21oi_1 _08934_ (.A1(_04086_),
    .A2(_04089_),
    .B1(_04085_),
    .Y(_04092_));
 sky130_fd_sc_hd__xor2_1 _08935_ (.A(_04091_),
    .B(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__nor2_1 _08936_ (.A(_04042_),
    .B(_04093_),
    .Y(net109));
 sky130_fd_sc_hd__or2_1 _08937_ (.A(_01384_),
    .B(\u_decod.branch_imm_q_o[18] ),
    .X(_04094_));
 sky130_fd_sc_hd__nand2_1 _08938_ (.A(_01384_),
    .B(\u_decod.branch_imm_q_o[18] ),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_1 _08939_ (.A(_04094_),
    .B(_04095_),
    .Y(_04096_));
 sky130_fd_sc_hd__o211a_1 _08940_ (.A1(_01380_),
    .A2(\u_decod.branch_imm_q_o[17] ),
    .B1(\u_decod.branch_imm_q_o[16] ),
    .C1(_01388_),
    .X(_04097_));
 sky130_fd_sc_hd__a21o_1 _08941_ (.A1(_01380_),
    .A2(\u_decod.branch_imm_q_o[17] ),
    .B1(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__a31oi_2 _08942_ (.A1(_04086_),
    .A2(_04089_),
    .A3(_04091_),
    .B1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__xnor2_1 _08943_ (.A(_04096_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__nor2_1 _08944_ (.A(_04042_),
    .B(_04100_),
    .Y(net110));
 sky130_fd_sc_hd__buf_2 _08945_ (.A(_02621_),
    .X(_04101_));
 sky130_fd_sc_hd__xor2_1 _08946_ (.A(_01376_),
    .B(\u_decod.branch_imm_q_o[19] ),
    .X(_04102_));
 sky130_fd_sc_hd__inv_2 _08947_ (.A(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__o21a_1 _08948_ (.A1(_04096_),
    .A2(_04099_),
    .B1(_04095_),
    .X(_04104_));
 sky130_fd_sc_hd__xnor2_1 _08949_ (.A(_04103_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__nor2_1 _08950_ (.A(_04101_),
    .B(_04105_),
    .Y(net111));
 sky130_fd_sc_hd__nand2_1 _08951_ (.A(_01363_),
    .B(\u_decod.branch_imm_q_o[20] ),
    .Y(_04106_));
 sky130_fd_sc_hd__or2_1 _08952_ (.A(_01363_),
    .B(\u_decod.branch_imm_q_o[20] ),
    .X(_04107_));
 sky130_fd_sc_hd__nand2_1 _08953_ (.A(_04106_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__o211a_1 _08954_ (.A1(_01376_),
    .A2(\u_decod.branch_imm_q_o[19] ),
    .B1(\u_decod.branch_imm_q_o[18] ),
    .C1(_01384_),
    .X(_04109_));
 sky130_fd_sc_hd__a21oi_1 _08955_ (.A1(_01376_),
    .A2(\u_decod.branch_imm_q_o[19] ),
    .B1(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__o31a_1 _08956_ (.A1(_04096_),
    .A2(_04099_),
    .A3(_04103_),
    .B1(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__xnor2_1 _08957_ (.A(_04108_),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _08958_ (.A(_04101_),
    .B(_04112_),
    .Y(net113));
 sky130_fd_sc_hd__xor2_1 _08959_ (.A(_01358_),
    .B(\u_decod.branch_imm_q_o[21] ),
    .X(_04113_));
 sky130_fd_sc_hd__inv_2 _08960_ (.A(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__o21a_1 _08961_ (.A1(_04108_),
    .A2(_04111_),
    .B1(_04106_),
    .X(_04115_));
 sky130_fd_sc_hd__xnor2_1 _08962_ (.A(_04114_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nor2_1 _08963_ (.A(_04101_),
    .B(_04116_),
    .Y(net114));
 sky130_fd_sc_hd__nand2_1 _08964_ (.A(_01371_),
    .B(\u_decod.branch_imm_q_o[22] ),
    .Y(_04117_));
 sky130_fd_sc_hd__or2_1 _08965_ (.A(_01371_),
    .B(\u_decod.branch_imm_q_o[22] ),
    .X(_04118_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_04117_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__o211a_1 _08967_ (.A1(_01358_),
    .A2(\u_decod.branch_imm_q_o[21] ),
    .B1(\u_decod.branch_imm_q_o[20] ),
    .C1(_01363_),
    .X(_04120_));
 sky130_fd_sc_hd__a21oi_1 _08968_ (.A1(_01358_),
    .A2(\u_decod.branch_imm_q_o[21] ),
    .B1(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__o31a_1 _08969_ (.A1(_04108_),
    .A2(_04111_),
    .A3(_04114_),
    .B1(_04121_),
    .X(_04122_));
 sky130_fd_sc_hd__xnor2_1 _08970_ (.A(_04119_),
    .B(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__nor2_1 _08971_ (.A(_04101_),
    .B(_04123_),
    .Y(net115));
 sky130_fd_sc_hd__or2_1 _08972_ (.A(_01367_),
    .B(\u_decod.branch_imm_q_o[23] ),
    .X(_04124_));
 sky130_fd_sc_hd__nand2_1 _08973_ (.A(_01367_),
    .B(\u_decod.branch_imm_q_o[23] ),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_04124_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__o21a_1 _08975_ (.A1(_04119_),
    .A2(_04122_),
    .B1(_04117_),
    .X(_04127_));
 sky130_fd_sc_hd__xnor2_1 _08976_ (.A(_04126_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__nor2_1 _08977_ (.A(_04101_),
    .B(_04128_),
    .Y(net116));
 sky130_fd_sc_hd__or2_1 _08978_ (.A(\u_decod.rs1_data_q[24] ),
    .B(\u_decod.branch_imm_q_o[24] ),
    .X(_04129_));
 sky130_fd_sc_hd__nand2_1 _08979_ (.A(\u_decod.rs1_data_q[24] ),
    .B(\u_decod.branch_imm_q_o[24] ),
    .Y(_04130_));
 sky130_fd_sc_hd__and2_1 _08980_ (.A(_04129_),
    .B(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__inv_2 _08981_ (.A(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__and3_1 _08982_ (.A(_01371_),
    .B(\u_decod.branch_imm_q_o[22] ),
    .C(_04124_),
    .X(_04133_));
 sky130_fd_sc_hd__a21oi_1 _08983_ (.A1(_01367_),
    .A2(\u_decod.branch_imm_q_o[23] ),
    .B1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__o31a_1 _08984_ (.A1(_04119_),
    .A2(_04122_),
    .A3(_04126_),
    .B1(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__xnor2_1 _08985_ (.A(_04132_),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_1 _08986_ (.A(_04101_),
    .B(_04136_),
    .Y(net117));
 sky130_fd_sc_hd__and2_1 _08987_ (.A(\u_decod.rs1_data_q[25] ),
    .B(\u_decod.branch_imm_q_o[25] ),
    .X(_04137_));
 sky130_fd_sc_hd__nor2_1 _08988_ (.A(\u_decod.rs1_data_q[25] ),
    .B(\u_decod.branch_imm_q_o[25] ),
    .Y(_04138_));
 sky130_fd_sc_hd__or2_1 _08989_ (.A(_04137_),
    .B(_04138_),
    .X(_04139_));
 sky130_fd_sc_hd__o21a_1 _08990_ (.A1(_04132_),
    .A2(_04135_),
    .B1(_04130_),
    .X(_04140_));
 sky130_fd_sc_hd__xnor2_1 _08991_ (.A(_04139_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__nor2_1 _08992_ (.A(_04101_),
    .B(_04141_),
    .Y(net118));
 sky130_fd_sc_hd__nand2_1 _08993_ (.A(\u_decod.rs1_data_q[26] ),
    .B(\u_decod.branch_imm_q_o[26] ),
    .Y(_04142_));
 sky130_fd_sc_hd__or2_1 _08994_ (.A(\u_decod.rs1_data_q[26] ),
    .B(\u_decod.branch_imm_q_o[26] ),
    .X(_04143_));
 sky130_fd_sc_hd__nand2_1 _08995_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__o21bai_1 _08996_ (.A1(_04138_),
    .A2(_04140_),
    .B1_N(_04137_),
    .Y(_04145_));
 sky130_fd_sc_hd__xor2_1 _08997_ (.A(_04144_),
    .B(_04145_),
    .X(_04146_));
 sky130_fd_sc_hd__nor2_1 _08998_ (.A(_04101_),
    .B(_04146_),
    .Y(net119));
 sky130_fd_sc_hd__or2_1 _08999_ (.A(\u_decod.rs1_data_q[27] ),
    .B(\u_decod.branch_imm_q_o[27] ),
    .X(_04147_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(\u_decod.rs1_data_q[27] ),
    .B(\u_decod.branch_imm_q_o[27] ),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(_04147_),
    .B(_04148_),
    .Y(_04149_));
 sky130_fd_sc_hd__a21bo_1 _09002_ (.A1(_04143_),
    .A2(_04145_),
    .B1_N(_04142_),
    .X(_04150_));
 sky130_fd_sc_hd__xor2_1 _09003_ (.A(_04149_),
    .B(_04150_),
    .X(_04151_));
 sky130_fd_sc_hd__nor2_1 _09004_ (.A(_04101_),
    .B(_04151_),
    .Y(net120));
 sky130_fd_sc_hd__or4_1 _09005_ (.A(_04132_),
    .B(_04139_),
    .C(_04144_),
    .D(_04149_),
    .X(_04152_));
 sky130_fd_sc_hd__a21oi_1 _09006_ (.A1(\u_decod.rs1_data_q[24] ),
    .A2(\u_decod.branch_imm_q_o[24] ),
    .B1(_04137_),
    .Y(_04153_));
 sky130_fd_sc_hd__a21bo_1 _09007_ (.A1(_04142_),
    .A2(_04148_),
    .B1_N(_04147_),
    .X(_04154_));
 sky130_fd_sc_hd__o41a_1 _09008_ (.A1(_04138_),
    .A2(_04144_),
    .A3(_04153_),
    .A4(_04149_),
    .B1(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__o21a_1 _09009_ (.A1(_04135_),
    .A2(_04152_),
    .B1(_04155_),
    .X(_04156_));
 sky130_fd_sc_hd__nor2_1 _09010_ (.A(\u_decod.rs1_data_q[28] ),
    .B(\u_decod.branch_imm_q_o[28] ),
    .Y(_04157_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(\u_decod.rs1_data_q[28] ),
    .B(\u_decod.branch_imm_q_o[28] ),
    .Y(_04158_));
 sky130_fd_sc_hd__and2b_1 _09012_ (.A_N(_04157_),
    .B(_04158_),
    .X(_04159_));
 sky130_fd_sc_hd__xor2_1 _09013_ (.A(_04156_),
    .B(_04159_),
    .X(_04160_));
 sky130_fd_sc_hd__nor2_1 _09014_ (.A(_04101_),
    .B(_04160_),
    .Y(net121));
 sky130_fd_sc_hd__or2_1 _09015_ (.A(\u_decod.rs1_data_q[29] ),
    .B(\u_decod.branch_imm_q_o[29] ),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(\u_decod.rs1_data_q[29] ),
    .B(\u_decod.branch_imm_q_o[29] ),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_1 _09017_ (.A(_04161_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__o21ai_1 _09018_ (.A1(_04156_),
    .A2(_04157_),
    .B1(_04158_),
    .Y(_04164_));
 sky130_fd_sc_hd__xor2_1 _09019_ (.A(_04163_),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__nor2_1 _09020_ (.A(_02621_),
    .B(_04165_),
    .Y(net122));
 sky130_fd_sc_hd__nand2_1 _09021_ (.A(\u_decod.rs1_data_q[30] ),
    .B(\u_decod.branch_imm_q_o[30] ),
    .Y(_04166_));
 sky130_fd_sc_hd__or2_1 _09022_ (.A(\u_decod.rs1_data_q[30] ),
    .B(\u_decod.branch_imm_q_o[30] ),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_1 _09023_ (.A(_04166_),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__a21boi_1 _09024_ (.A1(_04161_),
    .A2(_04164_),
    .B1_N(_04162_),
    .Y(_04169_));
 sky130_fd_sc_hd__xor2_1 _09025_ (.A(_04168_),
    .B(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__and2_1 _09026_ (.A(net133),
    .B(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__buf_1 _09027_ (.A(_04171_),
    .X(net124));
 sky130_fd_sc_hd__o21a_1 _09028_ (.A1(_04168_),
    .A2(_04169_),
    .B1(_04166_),
    .X(_04172_));
 sky130_fd_sc_hd__xor2_1 _09029_ (.A(_01267_),
    .B(\u_decod.branch_imm_q_o[31] ),
    .X(_04173_));
 sky130_fd_sc_hd__xnor2_1 _09030_ (.A(_04172_),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__and2_1 _09031_ (.A(net133),
    .B(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__buf_1 _09032_ (.A(_04175_),
    .X(net125));
 sky130_fd_sc_hd__and2_1 _09033_ (.A(_01420_),
    .B(_01421_),
    .X(_04176_));
 sky130_fd_sc_hd__or4b_1 _09034_ (.A(_01340_),
    .B(_01330_),
    .C(_01337_),
    .D_N(_01419_),
    .X(_04177_));
 sky130_fd_sc_hd__a211o_1 _09035_ (.A1(_01314_),
    .A2(_01426_),
    .B1(_01766_),
    .C1(_01813_),
    .X(_04178_));
 sky130_fd_sc_hd__or4_1 _09036_ (.A(_01350_),
    .B(_01345_),
    .C(_01342_),
    .D(_01347_),
    .X(_04179_));
 sky130_fd_sc_hd__or4_1 _09037_ (.A(_01355_),
    .B(_01352_),
    .C(_02588_),
    .D(_01391_),
    .X(_04180_));
 sky130_fd_sc_hd__nand4_1 _09038_ (.A(_01366_),
    .B(_01370_),
    .C(_01383_),
    .D(_01387_),
    .Y(_04181_));
 sky130_fd_sc_hd__or4b_1 _09039_ (.A(_01280_),
    .B(_01283_),
    .C(_01361_),
    .D_N(_01374_),
    .X(_04182_));
 sky130_fd_sc_hd__or4_1 _09040_ (.A(_04179_),
    .B(_04180_),
    .C(_04181_),
    .D(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__or4_1 _09041_ (.A(_01266_),
    .B(_01273_),
    .C(_01277_),
    .D(_01286_),
    .X(_04184_));
 sky130_fd_sc_hd__or4_2 _09042_ (.A(_01263_),
    .B(_01270_),
    .C(_04183_),
    .D(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__o211a_1 _09043_ (.A1(_01325_),
    .A2(_01326_),
    .B1(_01311_),
    .C1(_01316_),
    .X(_04186_));
 sky130_fd_sc_hd__or4b_1 _09044_ (.A(_01324_),
    .B(_04178_),
    .C(_04185_),
    .D_N(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__nor2_1 _09045_ (.A(_04177_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _09046_ (.A(\u_decod.unsign_ext_q_o ),
    .B(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__a21boi_1 _09047_ (.A1(_04176_),
    .A2(_04189_),
    .B1_N(\u_decod.instr_operation_q[3] ),
    .Y(_04190_));
 sky130_fd_sc_hd__o21a_1 _09048_ (.A1(_04177_),
    .A2(_04187_),
    .B1(_02781_),
    .X(_04191_));
 sky130_fd_sc_hd__a211o_1 _09049_ (.A1(\u_decod.instr_operation_q[0] ),
    .A2(_04188_),
    .B1(\u_decod.instr_operation_q[5] ),
    .C1(\u_decod.instr_operation_q[4] ),
    .X(_04192_));
 sky130_fd_sc_hd__a211o_1 _09050_ (.A1(_01430_),
    .A2(_04176_),
    .B1(_04191_),
    .C1(_04192_),
    .X(_04193_));
 sky130_fd_sc_hd__o21a_1 _09051_ (.A1(_04190_),
    .A2(_04193_),
    .B1(_01485_),
    .X(\u_exe.branch_v ));
 sky130_fd_sc_hd__inv_2 _09052_ (.A(\u_decod.instr_operation_q[5] ),
    .Y(_04194_));
 sky130_fd_sc_hd__and2_1 _09053_ (.A(_04194_),
    .B(\u_exe.branch_v ),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_2 _09054_ (.A(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_4 _09055_ (.A(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__nand2_1 _09056_ (.A(\u_decod.branch_imm_q_o[0] ),
    .B(\u_decod.pc_q_o[0] ),
    .Y(_04198_));
 sky130_fd_sc_hd__or2_1 _09057_ (.A(\u_decod.branch_imm_q_o[0] ),
    .B(\u_decod.pc_q_o[0] ),
    .X(_04199_));
 sky130_fd_sc_hd__nor2_2 _09058_ (.A(_04194_),
    .B(_02334_),
    .Y(_04200_));
 sky130_fd_sc_hd__inv_2 _09059_ (.A(_01066_),
    .Y(_04201_));
 sky130_fd_sc_hd__a32o_1 _09060_ (.A1(_04197_),
    .A2(_04198_),
    .A3(_04199_),
    .B1(_04200_),
    .B2(_04201_),
    .X(\u_exe.bu_pc_res[0] ));
 sky130_fd_sc_hd__nor2_1 _09061_ (.A(\u_decod.branch_imm_q_o[1] ),
    .B(\u_decod.pc_q_o[1] ),
    .Y(_04202_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(\u_decod.branch_imm_q_o[1] ),
    .B(\u_decod.pc_q_o[1] ),
    .Y(_04203_));
 sky130_fd_sc_hd__and2b_1 _09063_ (.A_N(_04202_),
    .B(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__xnor2_1 _09064_ (.A(_04198_),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__a22o_1 _09065_ (.A1(_01063_),
    .A2(_04200_),
    .B1(_04197_),
    .B2(_04205_),
    .X(\u_exe.bu_pc_res[1] ));
 sky130_fd_sc_hd__nand2_4 _09066_ (.A(\u_decod.instr_operation_q[5] ),
    .B(_01485_),
    .Y(_04206_));
 sky130_fd_sc_hd__buf_2 _09067_ (.A(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__buf_2 _09068_ (.A(_04196_),
    .X(_04208_));
 sky130_fd_sc_hd__o21a_1 _09069_ (.A1(_04198_),
    .A2(_04202_),
    .B1(_04203_),
    .X(_04209_));
 sky130_fd_sc_hd__nor2_1 _09070_ (.A(\u_decod.pc_q_o[2] ),
    .B(\u_decod.branch_imm_q_o[2] ),
    .Y(_04210_));
 sky130_fd_sc_hd__nand2_1 _09071_ (.A(\u_decod.pc_q_o[2] ),
    .B(\u_decod.branch_imm_q_o[2] ),
    .Y(_04211_));
 sky130_fd_sc_hd__and2b_1 _09072_ (.A_N(_04210_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__xnor2_1 _09073_ (.A(_04209_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__a2bb2o_1 _09074_ (.A1_N(_04004_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04213_),
    .X(\u_exe.bu_pc_res[2] ));
 sky130_fd_sc_hd__o211a_1 _09075_ (.A1(_04198_),
    .A2(_04202_),
    .B1(_04203_),
    .C1(_04211_),
    .X(_04214_));
 sky130_fd_sc_hd__nor2_1 _09076_ (.A(\u_decod.pc_q_o[3] ),
    .B(\u_decod.branch_imm_q_o[3] ),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _09077_ (.A(\u_decod.pc_q_o[3] ),
    .B(\u_decod.branch_imm_q_o[3] ),
    .Y(_04216_));
 sky130_fd_sc_hd__or2b_1 _09078_ (.A(_04215_),
    .B_N(_04216_),
    .X(_04217_));
 sky130_fd_sc_hd__o21ai_1 _09079_ (.A1(_04210_),
    .A2(_04214_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__or3_1 _09080_ (.A(_04210_),
    .B(_04217_),
    .C(_04214_),
    .X(_04219_));
 sky130_fd_sc_hd__nor2_1 _09081_ (.A(_04011_),
    .B(_04206_),
    .Y(_04220_));
 sky130_fd_sc_hd__a31o_1 _09082_ (.A1(_04197_),
    .A2(_04218_),
    .A3(_04219_),
    .B1(_04220_),
    .X(\u_exe.bu_pc_res[3] ));
 sky130_fd_sc_hd__nand2_1 _09083_ (.A(\u_decod.pc_q_o[4] ),
    .B(\u_decod.branch_imm_q_o[4] ),
    .Y(_04221_));
 sky130_fd_sc_hd__or2_1 _09084_ (.A(\u_decod.pc_q_o[4] ),
    .B(\u_decod.branch_imm_q_o[4] ),
    .X(_04222_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__o31a_1 _09086_ (.A1(_04210_),
    .A2(_04215_),
    .A3(_04214_),
    .B1(_04216_),
    .X(_04224_));
 sky130_fd_sc_hd__xor2_1 _09087_ (.A(_04223_),
    .B(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__a2bb2o_1 _09088_ (.A1_N(_04017_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04225_),
    .X(\u_exe.bu_pc_res[4] ));
 sky130_fd_sc_hd__nor2_1 _09089_ (.A(\u_decod.pc_q_o[5] ),
    .B(\u_decod.branch_imm_q_o[5] ),
    .Y(_04226_));
 sky130_fd_sc_hd__and2_1 _09090_ (.A(\u_decod.pc_q_o[5] ),
    .B(\u_decod.branch_imm_q_o[5] ),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_1 _09091_ (.A(_04226_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__o21a_1 _09092_ (.A1(_04223_),
    .A2(_04224_),
    .B1(_04221_),
    .X(_04229_));
 sky130_fd_sc_hd__xnor2_1 _09093_ (.A(_04228_),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__a2bb2o_1 _09094_ (.A1_N(_04022_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04230_),
    .X(\u_exe.bu_pc_res[5] ));
 sky130_fd_sc_hd__nand2_1 _09095_ (.A(\u_decod.pc_q_o[6] ),
    .B(\u_decod.branch_imm_q_o[6] ),
    .Y(_04231_));
 sky130_fd_sc_hd__or2_1 _09096_ (.A(\u_decod.pc_q_o[6] ),
    .B(\u_decod.branch_imm_q_o[6] ),
    .X(_04232_));
 sky130_fd_sc_hd__and2_1 _09097_ (.A(_04231_),
    .B(_04232_),
    .X(_04233_));
 sky130_fd_sc_hd__inv_2 _09098_ (.A(_04227_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand3b_1 _09099_ (.A_N(_04226_),
    .B(\u_decod.branch_imm_q_o[4] ),
    .C(\u_decod.pc_q_o[4] ),
    .Y(_04235_));
 sky130_fd_sc_hd__o311a_1 _09100_ (.A1(_04223_),
    .A2(_04224_),
    .A3(_04226_),
    .B1(_04234_),
    .C1(_04235_),
    .X(_04236_));
 sky130_fd_sc_hd__xnor2_1 _09101_ (.A(_04233_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__a2bb2o_1 _09102_ (.A1_N(_04029_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04237_),
    .X(\u_exe.bu_pc_res[6] ));
 sky130_fd_sc_hd__nor2_1 _09103_ (.A(\u_decod.pc_q_o[7] ),
    .B(\u_decod.branch_imm_q_o[7] ),
    .Y(_04238_));
 sky130_fd_sc_hd__nand2_1 _09104_ (.A(\u_decod.pc_q_o[7] ),
    .B(\u_decod.branch_imm_q_o[7] ),
    .Y(_04239_));
 sky130_fd_sc_hd__and2b_1 _09105_ (.A_N(_04238_),
    .B(_04239_),
    .X(_04240_));
 sky130_fd_sc_hd__inv_2 _09106_ (.A(_04233_),
    .Y(_04241_));
 sky130_fd_sc_hd__o21a_1 _09107_ (.A1(_04241_),
    .A2(_04236_),
    .B1(_04231_),
    .X(_04242_));
 sky130_fd_sc_hd__xnor2_1 _09108_ (.A(_04240_),
    .B(_04242_),
    .Y(_04243_));
 sky130_fd_sc_hd__a2bb2o_1 _09109_ (.A1_N(_04034_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04243_),
    .X(\u_exe.bu_pc_res[7] ));
 sky130_fd_sc_hd__or2_1 _09110_ (.A(\u_decod.pc_q_o[8] ),
    .B(\u_decod.branch_imm_q_o[8] ),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _09111_ (.A(\u_decod.pc_q_o[8] ),
    .B(\u_decod.branch_imm_q_o[8] ),
    .Y(_04245_));
 sky130_fd_sc_hd__and2_1 _09112_ (.A(_04244_),
    .B(_04245_),
    .X(_04246_));
 sky130_fd_sc_hd__nand3b_1 _09113_ (.A_N(_04238_),
    .B(\u_decod.branch_imm_q_o[6] ),
    .C(\u_decod.pc_q_o[6] ),
    .Y(_04247_));
 sky130_fd_sc_hd__o311a_1 _09114_ (.A1(_04241_),
    .A2(_04236_),
    .A3(_04238_),
    .B1(_04239_),
    .C1(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__xnor2_1 _09115_ (.A(_04246_),
    .B(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__a2bb2o_1 _09116_ (.A1_N(_04041_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04249_),
    .X(\u_exe.bu_pc_res[8] ));
 sky130_fd_sc_hd__nor2_1 _09117_ (.A(\u_decod.pc_q_o[9] ),
    .B(\u_decod.branch_imm_q_o[9] ),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _09118_ (.A(\u_decod.pc_q_o[9] ),
    .B(\u_decod.branch_imm_q_o[9] ),
    .Y(_04251_));
 sky130_fd_sc_hd__and2b_1 _09119_ (.A_N(_04250_),
    .B(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__inv_2 _09120_ (.A(_04246_),
    .Y(_04253_));
 sky130_fd_sc_hd__o21a_1 _09121_ (.A1(_04253_),
    .A2(_04248_),
    .B1(_04245_),
    .X(_04254_));
 sky130_fd_sc_hd__xnor2_1 _09122_ (.A(_04252_),
    .B(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__a2bb2o_1 _09123_ (.A1_N(_04047_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04255_),
    .X(\u_exe.bu_pc_res[9] ));
 sky130_fd_sc_hd__or2_1 _09124_ (.A(\u_decod.pc_q_o[10] ),
    .B(\u_decod.branch_imm_q_o[10] ),
    .X(_04256_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(\u_decod.pc_q_o[10] ),
    .B(\u_decod.branch_imm_q_o[10] ),
    .Y(_04257_));
 sky130_fd_sc_hd__and2_1 _09126_ (.A(_04256_),
    .B(_04257_),
    .X(_04258_));
 sky130_fd_sc_hd__nand3b_1 _09127_ (.A_N(_04250_),
    .B(\u_decod.branch_imm_q_o[8] ),
    .C(\u_decod.pc_q_o[8] ),
    .Y(_04259_));
 sky130_fd_sc_hd__o311a_1 _09128_ (.A1(_04253_),
    .A2(_04248_),
    .A3(_04250_),
    .B1(_04251_),
    .C1(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__xnor2_1 _09129_ (.A(_04258_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__a2bb2o_1 _09130_ (.A1_N(_04054_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04261_),
    .X(\u_exe.bu_pc_res[10] ));
 sky130_fd_sc_hd__nor2_1 _09131_ (.A(\u_decod.pc_q_o[11] ),
    .B(\u_decod.branch_imm_q_o[11] ),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(\u_decod.pc_q_o[11] ),
    .B(\u_decod.branch_imm_q_o[11] ),
    .Y(_04263_));
 sky130_fd_sc_hd__and2b_1 _09133_ (.A_N(_04262_),
    .B(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__inv_2 _09134_ (.A(_04258_),
    .Y(_04265_));
 sky130_fd_sc_hd__o21a_1 _09135_ (.A1(_04265_),
    .A2(_04260_),
    .B1(_04257_),
    .X(_04266_));
 sky130_fd_sc_hd__xnor2_1 _09136_ (.A(_04264_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a2bb2o_1 _09137_ (.A1_N(_04059_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04267_),
    .X(\u_exe.bu_pc_res[11] ));
 sky130_fd_sc_hd__or2_1 _09138_ (.A(\u_decod.pc_q_o[12] ),
    .B(\u_decod.branch_imm_q_o[12] ),
    .X(_04268_));
 sky130_fd_sc_hd__nand2_1 _09139_ (.A(\u_decod.pc_q_o[12] ),
    .B(\u_decod.branch_imm_q_o[12] ),
    .Y(_04269_));
 sky130_fd_sc_hd__and2_1 _09140_ (.A(_04268_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__nand3b_1 _09141_ (.A_N(_04262_),
    .B(\u_decod.branch_imm_q_o[10] ),
    .C(\u_decod.pc_q_o[10] ),
    .Y(_04271_));
 sky130_fd_sc_hd__o311a_1 _09142_ (.A1(_04265_),
    .A2(_04260_),
    .A3(_04262_),
    .B1(_04263_),
    .C1(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__xnor2_1 _09143_ (.A(_04270_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a2bb2o_1 _09144_ (.A1_N(_04066_),
    .A2_N(_04207_),
    .B1(_04208_),
    .B2(_04273_),
    .X(\u_exe.bu_pc_res[12] ));
 sky130_fd_sc_hd__clkbuf_2 _09145_ (.A(_04206_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_2 _09146_ (.A(_04196_),
    .X(_04275_));
 sky130_fd_sc_hd__nor2_1 _09147_ (.A(\u_decod.pc_q_o[13] ),
    .B(\u_decod.branch_imm_q_o[13] ),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(\u_decod.pc_q_o[13] ),
    .B(\u_decod.branch_imm_q_o[13] ),
    .Y(_04277_));
 sky130_fd_sc_hd__and2b_1 _09149_ (.A_N(_04276_),
    .B(_04277_),
    .X(_04278_));
 sky130_fd_sc_hd__inv_2 _09150_ (.A(_04270_),
    .Y(_04279_));
 sky130_fd_sc_hd__o21a_1 _09151_ (.A1(_04279_),
    .A2(_04272_),
    .B1(_04269_),
    .X(_04280_));
 sky130_fd_sc_hd__xnor2_1 _09152_ (.A(_04278_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__a2bb2o_1 _09153_ (.A1_N(_04071_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04281_),
    .X(\u_exe.bu_pc_res[13] ));
 sky130_fd_sc_hd__or2_1 _09154_ (.A(\u_decod.pc_q_o[14] ),
    .B(\u_decod.branch_imm_q_o[14] ),
    .X(_04282_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(\u_decod.pc_q_o[14] ),
    .B(\u_decod.branch_imm_q_o[14] ),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _09156_ (.A(_04282_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand3b_1 _09157_ (.A_N(_04276_),
    .B(\u_decod.branch_imm_q_o[12] ),
    .C(\u_decod.pc_q_o[12] ),
    .Y(_04285_));
 sky130_fd_sc_hd__o311a_1 _09158_ (.A1(_04279_),
    .A2(_04272_),
    .A3(_04276_),
    .B1(_04277_),
    .C1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__or2_1 _09159_ (.A(_04284_),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__nand2_1 _09160_ (.A(_04284_),
    .B(_04286_),
    .Y(_04288_));
 sky130_fd_sc_hd__and2_1 _09161_ (.A(_04287_),
    .B(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__a2bb2o_1 _09162_ (.A1_N(_04078_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04289_),
    .X(\u_exe.bu_pc_res[14] ));
 sky130_fd_sc_hd__nor2_1 _09163_ (.A(\u_decod.pc_q_o[15] ),
    .B(\u_decod.branch_imm_q_o[15] ),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(\u_decod.pc_q_o[15] ),
    .B(\u_decod.branch_imm_q_o[15] ),
    .Y(_04291_));
 sky130_fd_sc_hd__and2b_1 _09165_ (.A_N(_04290_),
    .B(_04291_),
    .X(_04292_));
 sky130_fd_sc_hd__and2_1 _09166_ (.A(_04283_),
    .B(_04287_),
    .X(_04293_));
 sky130_fd_sc_hd__xnor2_1 _09167_ (.A(_04292_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__a2bb2o_1 _09168_ (.A1_N(_04083_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04294_),
    .X(\u_exe.bu_pc_res[15] ));
 sky130_fd_sc_hd__or2_1 _09169_ (.A(\u_decod.pc_q_o[16] ),
    .B(\u_decod.branch_imm_q_o[16] ),
    .X(_04295_));
 sky130_fd_sc_hd__nand2_1 _09170_ (.A(\u_decod.pc_q_o[16] ),
    .B(\u_decod.branch_imm_q_o[16] ),
    .Y(_04296_));
 sky130_fd_sc_hd__nand2_1 _09171_ (.A(_04295_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__a31o_1 _09172_ (.A1(_04283_),
    .A2(_04287_),
    .A3(_04291_),
    .B1(_04290_),
    .X(_04298_));
 sky130_fd_sc_hd__xor2_1 _09173_ (.A(_04297_),
    .B(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__a2bb2o_1 _09174_ (.A1_N(_04090_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04299_),
    .X(\u_exe.bu_pc_res[16] ));
 sky130_fd_sc_hd__nor2_1 _09175_ (.A(\u_decod.pc_q_o[17] ),
    .B(\u_decod.branch_imm_q_o[17] ),
    .Y(_04300_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(\u_decod.pc_q_o[17] ),
    .B(\u_decod.branch_imm_q_o[17] ),
    .Y(_04301_));
 sky130_fd_sc_hd__or2b_1 _09177_ (.A(_04300_),
    .B_N(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__a311o_1 _09178_ (.A1(_04283_),
    .A2(_04287_),
    .A3(_04291_),
    .B1(_04297_),
    .C1(_04290_),
    .X(_04303_));
 sky130_fd_sc_hd__nand2_1 _09179_ (.A(_04296_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__xnor2_1 _09180_ (.A(_04302_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__a2bb2o_1 _09181_ (.A1_N(_04093_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04305_),
    .X(\u_exe.bu_pc_res[17] ));
 sky130_fd_sc_hd__or2_1 _09182_ (.A(\u_decod.pc_q_o[18] ),
    .B(\u_decod.branch_imm_q_o[18] ),
    .X(_04306_));
 sky130_fd_sc_hd__nand2_1 _09183_ (.A(\u_decod.pc_q_o[18] ),
    .B(\u_decod.branch_imm_q_o[18] ),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(_04306_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__a31o_1 _09185_ (.A1(_04296_),
    .A2(_04303_),
    .A3(_04301_),
    .B1(_04300_),
    .X(_04309_));
 sky130_fd_sc_hd__xor2_1 _09186_ (.A(_04308_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__a2bb2o_1 _09187_ (.A1_N(_04100_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04310_),
    .X(\u_exe.bu_pc_res[18] ));
 sky130_fd_sc_hd__nor2_1 _09188_ (.A(\u_decod.pc_q_o[19] ),
    .B(\u_decod.branch_imm_q_o[19] ),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _09189_ (.A(\u_decod.pc_q_o[19] ),
    .B(\u_decod.branch_imm_q_o[19] ),
    .Y(_04312_));
 sky130_fd_sc_hd__or2b_1 _09190_ (.A(_04311_),
    .B_N(_04312_),
    .X(_04313_));
 sky130_fd_sc_hd__a311o_1 _09191_ (.A1(_04296_),
    .A2(_04303_),
    .A3(_04301_),
    .B1(_04308_),
    .C1(_04300_),
    .X(_04314_));
 sky130_fd_sc_hd__nand2_1 _09192_ (.A(_04307_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__xnor2_1 _09193_ (.A(_04313_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__a2bb2o_1 _09194_ (.A1_N(_04105_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04316_),
    .X(\u_exe.bu_pc_res[19] ));
 sky130_fd_sc_hd__or2_1 _09195_ (.A(\u_decod.pc_q_o[20] ),
    .B(\u_decod.branch_imm_q_o[20] ),
    .X(_04317_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(\u_decod.pc_q_o[20] ),
    .B(\u_decod.branch_imm_q_o[20] ),
    .Y(_04318_));
 sky130_fd_sc_hd__nand2_1 _09197_ (.A(_04317_),
    .B(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__a311o_1 _09198_ (.A1(_04307_),
    .A2(_04314_),
    .A3(_04312_),
    .B1(_04319_),
    .C1(_04311_),
    .X(_04320_));
 sky130_fd_sc_hd__a31o_1 _09199_ (.A1(_04307_),
    .A2(_04314_),
    .A3(_04312_),
    .B1(_04311_),
    .X(_04321_));
 sky130_fd_sc_hd__a21boi_1 _09200_ (.A1(_04319_),
    .A2(_04321_),
    .B1_N(_04196_),
    .Y(_04322_));
 sky130_fd_sc_hd__a2bb2o_1 _09201_ (.A1_N(_04112_),
    .A2_N(_04274_),
    .B1(_04320_),
    .B2(_04322_),
    .X(\u_exe.bu_pc_res[20] ));
 sky130_fd_sc_hd__nor2_1 _09202_ (.A(\u_decod.pc_q_o[21] ),
    .B(\u_decod.branch_imm_q_o[21] ),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(\u_decod.pc_q_o[21] ),
    .B(\u_decod.branch_imm_q_o[21] ),
    .Y(_04324_));
 sky130_fd_sc_hd__or2b_1 _09204_ (.A(_04323_),
    .B_N(_04324_),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _09205_ (.A(_04318_),
    .B(_04320_),
    .Y(_04326_));
 sky130_fd_sc_hd__xnor2_1 _09206_ (.A(_04325_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__a2bb2o_1 _09207_ (.A1_N(_04116_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04327_),
    .X(\u_exe.bu_pc_res[21] ));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(\u_decod.pc_q_o[22] ),
    .B(\u_decod.branch_imm_q_o[22] ),
    .Y(_04328_));
 sky130_fd_sc_hd__or2_1 _09209_ (.A(\u_decod.pc_q_o[22] ),
    .B(\u_decod.branch_imm_q_o[22] ),
    .X(_04329_));
 sky130_fd_sc_hd__nand2_1 _09210_ (.A(_04328_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a311o_1 _09211_ (.A1(_04318_),
    .A2(_04320_),
    .A3(_04324_),
    .B1(_04330_),
    .C1(_04323_),
    .X(_04331_));
 sky130_fd_sc_hd__a31o_1 _09212_ (.A1(_04318_),
    .A2(_04320_),
    .A3(_04324_),
    .B1(_04323_),
    .X(_04332_));
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(_04330_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__nor2_1 _09214_ (.A(_04123_),
    .B(_04206_),
    .Y(_04334_));
 sky130_fd_sc_hd__a31o_1 _09215_ (.A1(_04197_),
    .A2(_04331_),
    .A3(_04333_),
    .B1(_04334_),
    .X(\u_exe.bu_pc_res[22] ));
 sky130_fd_sc_hd__nor2_1 _09216_ (.A(\u_decod.pc_q_o[23] ),
    .B(\u_decod.branch_imm_q_o[23] ),
    .Y(_04335_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(\u_decod.pc_q_o[23] ),
    .B(\u_decod.branch_imm_q_o[23] ),
    .Y(_04336_));
 sky130_fd_sc_hd__or2b_1 _09218_ (.A(_04335_),
    .B_N(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__nand2_1 _09219_ (.A(_04328_),
    .B(_04331_),
    .Y(_04338_));
 sky130_fd_sc_hd__xnor2_1 _09220_ (.A(_04337_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__a2bb2o_1 _09221_ (.A1_N(_04128_),
    .A2_N(_04274_),
    .B1(_04275_),
    .B2(_04339_),
    .X(\u_exe.bu_pc_res[23] ));
 sky130_fd_sc_hd__nand2_1 _09222_ (.A(\u_decod.pc_q_o[24] ),
    .B(\u_decod.branch_imm_q_o[24] ),
    .Y(_04340_));
 sky130_fd_sc_hd__or2_1 _09223_ (.A(\u_decod.pc_q_o[24] ),
    .B(\u_decod.branch_imm_q_o[24] ),
    .X(_04341_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(_04340_),
    .B(_04341_),
    .Y(_04342_));
 sky130_fd_sc_hd__a31o_1 _09225_ (.A1(_04328_),
    .A2(_04331_),
    .A3(_04336_),
    .B1(_04335_),
    .X(_04343_));
 sky130_fd_sc_hd__xor2_1 _09226_ (.A(_04342_),
    .B(_04343_),
    .X(_04344_));
 sky130_fd_sc_hd__a2bb2o_1 _09227_ (.A1_N(_04136_),
    .A2_N(_04206_),
    .B1(_04275_),
    .B2(_04344_),
    .X(\u_exe.bu_pc_res[24] ));
 sky130_fd_sc_hd__nand2_1 _09228_ (.A(\u_decod.pc_q_o[25] ),
    .B(\u_decod.branch_imm_q_o[25] ),
    .Y(_04345_));
 sky130_fd_sc_hd__or2_1 _09229_ (.A(\u_decod.pc_q_o[25] ),
    .B(\u_decod.branch_imm_q_o[25] ),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__o21a_1 _09231_ (.A1(_04342_),
    .A2(_04343_),
    .B1(_04340_),
    .X(_04348_));
 sky130_fd_sc_hd__xor2_1 _09232_ (.A(_04347_),
    .B(_04348_),
    .X(_04349_));
 sky130_fd_sc_hd__a2bb2o_1 _09233_ (.A1_N(_04141_),
    .A2_N(_04206_),
    .B1(_04197_),
    .B2(_04349_),
    .X(\u_exe.bu_pc_res[25] ));
 sky130_fd_sc_hd__nand2_1 _09234_ (.A(\u_decod.pc_q_o[26] ),
    .B(\u_decod.branch_imm_q_o[26] ),
    .Y(_04350_));
 sky130_fd_sc_hd__or2_1 _09235_ (.A(\u_decod.pc_q_o[26] ),
    .B(\u_decod.branch_imm_q_o[26] ),
    .X(_04351_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_04350_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__a21boi_1 _09237_ (.A1(_04345_),
    .A2(_04348_),
    .B1_N(_04346_),
    .Y(_04353_));
 sky130_fd_sc_hd__xnor2_1 _09238_ (.A(_04352_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__a2bb2o_1 _09239_ (.A1_N(_04146_),
    .A2_N(_04206_),
    .B1(_04197_),
    .B2(_04354_),
    .X(\u_exe.bu_pc_res[26] ));
 sky130_fd_sc_hd__and2_1 _09240_ (.A(\u_decod.pc_q_o[27] ),
    .B(\u_decod.branch_imm_q_o[27] ),
    .X(_04355_));
 sky130_fd_sc_hd__nor2_1 _09241_ (.A(\u_decod.pc_q_o[27] ),
    .B(\u_decod.branch_imm_q_o[27] ),
    .Y(_04356_));
 sky130_fd_sc_hd__nor2_1 _09242_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__a21boi_1 _09243_ (.A1(_04351_),
    .A2(_04353_),
    .B1_N(_04350_),
    .Y(_04358_));
 sky130_fd_sc_hd__xnor2_1 _09244_ (.A(_04357_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__a2bb2o_1 _09245_ (.A1_N(_04151_),
    .A2_N(_04206_),
    .B1(_04197_),
    .B2(_04359_),
    .X(\u_exe.bu_pc_res[27] ));
 sky130_fd_sc_hd__or3_1 _09246_ (.A(_04352_),
    .B(_04355_),
    .C(_04356_),
    .X(_04360_));
 sky130_fd_sc_hd__or3_1 _09247_ (.A(_04342_),
    .B(_04347_),
    .C(_04360_),
    .X(_04361_));
 sky130_fd_sc_hd__a311o_1 _09248_ (.A1(_04328_),
    .A2(_04331_),
    .A3(_04336_),
    .B1(_04361_),
    .C1(_04335_),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _09249_ (.A(_04340_),
    .B(_04345_),
    .Y(_04363_));
 sky130_fd_sc_hd__and3b_1 _09250_ (.A_N(_04360_),
    .B(_04363_),
    .C(_04346_),
    .X(_04364_));
 sky130_fd_sc_hd__inv_2 _09251_ (.A(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__o21ba_1 _09252_ (.A1(_04350_),
    .A2(_04356_),
    .B1_N(_04355_),
    .X(_04366_));
 sky130_fd_sc_hd__nand3_1 _09253_ (.A(_04362_),
    .B(_04365_),
    .C(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__nor2_1 _09254_ (.A(\u_decod.pc_q_o[28] ),
    .B(\u_decod.branch_imm_q_o[28] ),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(\u_decod.pc_q_o[28] ),
    .B(\u_decod.branch_imm_q_o[28] ),
    .Y(_04369_));
 sky130_fd_sc_hd__or2b_1 _09256_ (.A(_04368_),
    .B_N(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__xnor2_1 _09257_ (.A(_04367_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__a2bb2o_1 _09258_ (.A1_N(_04160_),
    .A2_N(_04206_),
    .B1(_04197_),
    .B2(_04371_),
    .X(\u_exe.bu_pc_res[28] ));
 sky130_fd_sc_hd__nor2_1 _09259_ (.A(\u_decod.pc_q_o[29] ),
    .B(\u_decod.branch_imm_q_o[29] ),
    .Y(_04372_));
 sky130_fd_sc_hd__and2_1 _09260_ (.A(\u_decod.pc_q_o[29] ),
    .B(\u_decod.branch_imm_q_o[29] ),
    .X(_04373_));
 sky130_fd_sc_hd__a41o_1 _09261_ (.A1(_04362_),
    .A2(_04365_),
    .A3(_04366_),
    .A4(_04369_),
    .B1(_04368_),
    .X(_04374_));
 sky130_fd_sc_hd__o21ai_1 _09262_ (.A1(_04372_),
    .A2(_04373_),
    .B1(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__o31a_1 _09263_ (.A1(_04372_),
    .A2(_04373_),
    .A3(_04374_),
    .B1(_04196_),
    .X(_04376_));
 sky130_fd_sc_hd__a2bb2o_1 _09264_ (.A1_N(_04165_),
    .A2_N(_04206_),
    .B1(_04375_),
    .B2(_04376_),
    .X(\u_exe.bu_pc_res[29] ));
 sky130_fd_sc_hd__or2_1 _09265_ (.A(\u_decod.pc_q_o[30] ),
    .B(\u_decod.branch_imm_q_o[30] ),
    .X(_04377_));
 sky130_fd_sc_hd__nand2_1 _09266_ (.A(\u_decod.pc_q_o[30] ),
    .B(\u_decod.branch_imm_q_o[30] ),
    .Y(_04378_));
 sky130_fd_sc_hd__nor2_1 _09267_ (.A(_04372_),
    .B(_04374_),
    .Y(_04379_));
 sky130_fd_sc_hd__a211o_1 _09268_ (.A1(_04377_),
    .A2(_04378_),
    .B1(_04379_),
    .C1(_04373_),
    .X(_04380_));
 sky130_fd_sc_hd__o211ai_2 _09269_ (.A1(_04373_),
    .A2(_04379_),
    .B1(_04378_),
    .C1(_04377_),
    .Y(_04381_));
 sky130_fd_sc_hd__a32o_1 _09270_ (.A1(_04197_),
    .A2(_04380_),
    .A3(_04381_),
    .B1(_04200_),
    .B2(_04170_),
    .X(\u_exe.bu_pc_res[30] ));
 sky130_fd_sc_hd__xnor2_1 _09271_ (.A(\u_decod.pc_q_o[31] ),
    .B(\u_decod.branch_imm_q_o[31] ),
    .Y(_04382_));
 sky130_fd_sc_hd__nand3_1 _09272_ (.A(_04378_),
    .B(_04381_),
    .C(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21o_1 _09273_ (.A1(_04378_),
    .A2(_04381_),
    .B1(_04382_),
    .X(_04384_));
 sky130_fd_sc_hd__a32o_1 _09274_ (.A1(_04197_),
    .A2(_04383_),
    .A3(_04384_),
    .B1(_04200_),
    .B2(_04174_),
    .X(\u_exe.bu_pc_res[31] ));
 sky130_fd_sc_hd__nor2_1 _09275_ (.A(_01481_),
    .B(_03998_),
    .Y(net167));
 sky130_fd_sc_hd__nor2_2 _09276_ (.A(_01477_),
    .B(_03998_),
    .Y(net178));
 sky130_fd_sc_hd__nor2_2 _09277_ (.A(_02685_),
    .B(_03998_),
    .Y(net189));
 sky130_fd_sc_hd__clkbuf_2 _09278_ (.A(\u_decod.instr_unit_q[3] ),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_2 _09279_ (.A(_01427_),
    .X(_04386_));
 sky130_fd_sc_hd__and3_1 _09280_ (.A(_04385_),
    .B(_01469_),
    .C(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__buf_1 _09281_ (.A(_04387_),
    .X(net192));
 sky130_fd_sc_hd__and3_1 _09282_ (.A(_04385_),
    .B(_01466_),
    .C(_04386_),
    .X(_04388_));
 sky130_fd_sc_hd__buf_1 _09283_ (.A(_04388_),
    .X(net193));
 sky130_fd_sc_hd__and3_1 _09284_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[5] ),
    .C(_04386_),
    .X(_04389_));
 sky130_fd_sc_hd__buf_1 _09285_ (.A(_04389_),
    .X(net194));
 sky130_fd_sc_hd__and3_1 _09286_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[6] ),
    .C(_04386_),
    .X(_04390_));
 sky130_fd_sc_hd__buf_1 _09287_ (.A(_04390_),
    .X(net195));
 sky130_fd_sc_hd__and3_1 _09288_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[7] ),
    .C(_04386_),
    .X(_04391_));
 sky130_fd_sc_hd__buf_1 _09289_ (.A(_04391_),
    .X(net196));
 sky130_fd_sc_hd__and3_1 _09290_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[8] ),
    .C(_04386_),
    .X(_04392_));
 sky130_fd_sc_hd__buf_1 _09291_ (.A(_04392_),
    .X(net197));
 sky130_fd_sc_hd__and3_1 _09292_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[9] ),
    .C(_04386_),
    .X(_04393_));
 sky130_fd_sc_hd__buf_1 _09293_ (.A(_04393_),
    .X(net198));
 sky130_fd_sc_hd__and3_1 _09294_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[10] ),
    .C(_04386_),
    .X(_04394_));
 sky130_fd_sc_hd__buf_1 _09295_ (.A(_04394_),
    .X(net168));
 sky130_fd_sc_hd__and3_1 _09296_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[11] ),
    .C(_04386_),
    .X(_04395_));
 sky130_fd_sc_hd__buf_1 _09297_ (.A(_04395_),
    .X(net169));
 sky130_fd_sc_hd__and3_1 _09298_ (.A(_04385_),
    .B(\u_decod.rs2_data_q[12] ),
    .C(_04386_),
    .X(_04396_));
 sky130_fd_sc_hd__buf_1 _09299_ (.A(_04396_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 _09300_ (.A(\u_decod.instr_unit_q[3] ),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_2 _09301_ (.A(_01427_),
    .X(_04398_));
 sky130_fd_sc_hd__and3_1 _09302_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[13] ),
    .C(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_2 _09303_ (.A(_04399_),
    .X(net171));
 sky130_fd_sc_hd__and3_1 _09304_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[14] ),
    .C(_04398_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_2 _09305_ (.A(_04400_),
    .X(net172));
 sky130_fd_sc_hd__and3_1 _09306_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[15] ),
    .C(_04398_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_2 _09307_ (.A(_04401_),
    .X(net173));
 sky130_fd_sc_hd__and3_1 _09308_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[16] ),
    .C(_04398_),
    .X(_04402_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09309_ (.A(_04402_),
    .X(net174));
 sky130_fd_sc_hd__and3_1 _09310_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[17] ),
    .C(_04398_),
    .X(_04403_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09311_ (.A(_04403_),
    .X(net175));
 sky130_fd_sc_hd__and3_1 _09312_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[18] ),
    .C(_04398_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_2 _09313_ (.A(_04404_),
    .X(net176));
 sky130_fd_sc_hd__and3_1 _09314_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[19] ),
    .C(_04398_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_2 _09315_ (.A(_04405_),
    .X(net177));
 sky130_fd_sc_hd__and3_1 _09316_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[20] ),
    .C(_04398_),
    .X(_04406_));
 sky130_fd_sc_hd__clkbuf_2 _09317_ (.A(_04406_),
    .X(net179));
 sky130_fd_sc_hd__and3_1 _09318_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[21] ),
    .C(_04398_),
    .X(_04407_));
 sky130_fd_sc_hd__clkbuf_2 _09319_ (.A(_04407_),
    .X(net180));
 sky130_fd_sc_hd__and3_1 _09320_ (.A(_04397_),
    .B(\u_decod.rs2_data_q[22] ),
    .C(_04398_),
    .X(_04408_));
 sky130_fd_sc_hd__clkbuf_2 _09321_ (.A(_04408_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 _09322_ (.A(\u_decod.instr_unit_q[3] ),
    .X(_04409_));
 sky130_fd_sc_hd__clkbuf_2 _09323_ (.A(_01427_),
    .X(_04410_));
 sky130_fd_sc_hd__and3_1 _09324_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[23] ),
    .C(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09325_ (.A(_04411_),
    .X(net182));
 sky130_fd_sc_hd__and3_1 _09326_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[24] ),
    .C(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__buf_1 _09327_ (.A(_04412_),
    .X(net183));
 sky130_fd_sc_hd__and3_1 _09328_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[25] ),
    .C(_04410_),
    .X(_04413_));
 sky130_fd_sc_hd__buf_1 _09329_ (.A(_04413_),
    .X(net184));
 sky130_fd_sc_hd__and3_1 _09330_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[26] ),
    .C(_04410_),
    .X(_04414_));
 sky130_fd_sc_hd__buf_1 _09331_ (.A(_04414_),
    .X(net185));
 sky130_fd_sc_hd__and3_1 _09332_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[27] ),
    .C(_04410_),
    .X(_04415_));
 sky130_fd_sc_hd__buf_1 _09333_ (.A(_04415_),
    .X(net186));
 sky130_fd_sc_hd__and3_1 _09334_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[28] ),
    .C(_04410_),
    .X(_04416_));
 sky130_fd_sc_hd__buf_1 _09335_ (.A(_04416_),
    .X(net187));
 sky130_fd_sc_hd__and3_1 _09336_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[29] ),
    .C(_04410_),
    .X(_04417_));
 sky130_fd_sc_hd__buf_1 _09337_ (.A(_04417_),
    .X(net188));
 sky130_fd_sc_hd__and3_1 _09338_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[30] ),
    .C(_04410_),
    .X(_04418_));
 sky130_fd_sc_hd__buf_1 _09339_ (.A(_04418_),
    .X(net190));
 sky130_fd_sc_hd__and3_1 _09340_ (.A(_04409_),
    .B(\u_decod.rs2_data_q[31] ),
    .C(_04410_),
    .X(_04419_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _09341_ (.A(_04419_),
    .X(net191));
 sky130_fd_sc_hd__and3_1 _09342_ (.A(_04409_),
    .B(\u_decod.instr_operation_q[0] ),
    .C(_04410_),
    .X(_04420_));
 sky130_fd_sc_hd__buf_1 _09343_ (.A(_04420_),
    .X(net166));
 sky130_fd_sc_hd__buf_2 _09344_ (.A(\u_decod.rf_ff_res_data_i[0] ),
    .X(_04421_));
 sky130_fd_sc_hd__nand2_1 _09345_ (.A(_01539_),
    .B(\u_decod.rf_write_v_q_i ),
    .Y(_04422_));
 sky130_fd_sc_hd__buf_4 _09346_ (.A(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__buf_2 _09347_ (.A(\u_decod.rf_ff_rd_adr_q_i[1] ),
    .X(_04424_));
 sky130_fd_sc_hd__nand2_1 _09348_ (.A(_01534_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__or3_2 _09349_ (.A(_01531_),
    .B(_01536_),
    .C(_04425_),
    .X(_04426_));
 sky130_fd_sc_hd__nor2_4 _09350_ (.A(_04423_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__clkbuf_8 _09351_ (.A(_04427_),
    .X(_04428_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(\u_rf.reg2_q[0] ),
    .A1(_04421_),
    .S(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _09353_ (.A(_04429_),
    .X(_00000_));
 sky130_fd_sc_hd__buf_2 _09354_ (.A(\u_decod.rf_ff_res_data_i[1] ),
    .X(_04430_));
 sky130_fd_sc_hd__mux2_1 _09355_ (.A0(\u_rf.reg2_q[1] ),
    .A1(_04430_),
    .S(_04428_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _09356_ (.A(_04431_),
    .X(_00001_));
 sky130_fd_sc_hd__buf_2 _09357_ (.A(\u_decod.rf_ff_res_data_i[2] ),
    .X(_04432_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(\u_rf.reg2_q[2] ),
    .A1(_04432_),
    .S(_04428_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _09359_ (.A(_04433_),
    .X(_00002_));
 sky130_fd_sc_hd__buf_2 _09360_ (.A(\u_decod.rf_ff_res_data_i[3] ),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _09361_ (.A0(\u_rf.reg2_q[3] ),
    .A1(_04434_),
    .S(_04428_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _09362_ (.A(_04435_),
    .X(_00003_));
 sky130_fd_sc_hd__buf_2 _09363_ (.A(\u_decod.rf_ff_res_data_i[4] ),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(\u_rf.reg2_q[4] ),
    .A1(_04436_),
    .S(_04428_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _09365_ (.A(_04437_),
    .X(_00004_));
 sky130_fd_sc_hd__buf_2 _09366_ (.A(\u_decod.rf_ff_res_data_i[5] ),
    .X(_04438_));
 sky130_fd_sc_hd__mux2_1 _09367_ (.A0(\u_rf.reg2_q[5] ),
    .A1(_04438_),
    .S(_04428_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _09368_ (.A(_04439_),
    .X(_00005_));
 sky130_fd_sc_hd__buf_2 _09369_ (.A(\u_decod.rf_ff_res_data_i[6] ),
    .X(_04440_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(\u_rf.reg2_q[6] ),
    .A1(_04440_),
    .S(_04428_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _09371_ (.A(_04441_),
    .X(_00006_));
 sky130_fd_sc_hd__clkbuf_2 _09372_ (.A(\u_decod.rf_ff_res_data_i[7] ),
    .X(_04442_));
 sky130_fd_sc_hd__mux2_1 _09373_ (.A0(\u_rf.reg2_q[7] ),
    .A1(_04442_),
    .S(_04428_),
    .X(_04443_));
 sky130_fd_sc_hd__clkbuf_1 _09374_ (.A(_04443_),
    .X(_00007_));
 sky130_fd_sc_hd__buf_2 _09375_ (.A(\u_decod.rf_ff_res_data_i[8] ),
    .X(_04444_));
 sky130_fd_sc_hd__mux2_1 _09376_ (.A0(\u_rf.reg2_q[8] ),
    .A1(_04444_),
    .S(_04428_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _09377_ (.A(_04445_),
    .X(_00008_));
 sky130_fd_sc_hd__buf_2 _09378_ (.A(\u_decod.rf_ff_res_data_i[9] ),
    .X(_04446_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(\u_rf.reg2_q[9] ),
    .A1(_04446_),
    .S(_04428_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _09380_ (.A(_04447_),
    .X(_00009_));
 sky130_fd_sc_hd__buf_2 _09381_ (.A(\u_decod.rf_ff_res_data_i[10] ),
    .X(_04448_));
 sky130_fd_sc_hd__buf_6 _09382_ (.A(_04427_),
    .X(_04449_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(\u_rf.reg2_q[10] ),
    .A1(_04448_),
    .S(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _09384_ (.A(_04450_),
    .X(_00010_));
 sky130_fd_sc_hd__clkbuf_2 _09385_ (.A(\u_decod.rf_ff_res_data_i[11] ),
    .X(_04451_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(\u_rf.reg2_q[11] ),
    .A1(_04451_),
    .S(_04449_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _09387_ (.A(_04452_),
    .X(_00011_));
 sky130_fd_sc_hd__clkbuf_2 _09388_ (.A(\u_decod.rf_ff_res_data_i[12] ),
    .X(_04453_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(\u_rf.reg2_q[12] ),
    .A1(_04453_),
    .S(_04449_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _09390_ (.A(_04454_),
    .X(_00012_));
 sky130_fd_sc_hd__clkbuf_2 _09391_ (.A(\u_decod.rf_ff_res_data_i[13] ),
    .X(_04455_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(\u_rf.reg2_q[13] ),
    .A1(_04455_),
    .S(_04449_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _09393_ (.A(_04456_),
    .X(_00013_));
 sky130_fd_sc_hd__buf_2 _09394_ (.A(\u_decod.rf_ff_res_data_i[14] ),
    .X(_04457_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(\u_rf.reg2_q[14] ),
    .A1(_04457_),
    .S(_04449_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _09396_ (.A(_04458_),
    .X(_00014_));
 sky130_fd_sc_hd__clkbuf_2 _09397_ (.A(\u_decod.rf_ff_res_data_i[15] ),
    .X(_04459_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(\u_rf.reg2_q[15] ),
    .A1(_04459_),
    .S(_04449_),
    .X(_04460_));
 sky130_fd_sc_hd__clkbuf_1 _09399_ (.A(_04460_),
    .X(_00015_));
 sky130_fd_sc_hd__buf_2 _09400_ (.A(\u_decod.rf_ff_res_data_i[16] ),
    .X(_04461_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(\u_rf.reg2_q[16] ),
    .A1(_04461_),
    .S(_04449_),
    .X(_04462_));
 sky130_fd_sc_hd__clkbuf_1 _09402_ (.A(_04462_),
    .X(_00016_));
 sky130_fd_sc_hd__buf_2 _09403_ (.A(\u_decod.rf_ff_res_data_i[17] ),
    .X(_04463_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(\u_rf.reg2_q[17] ),
    .A1(_04463_),
    .S(_04449_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _09405_ (.A(_04464_),
    .X(_00017_));
 sky130_fd_sc_hd__clkbuf_2 _09406_ (.A(\u_decod.rf_ff_res_data_i[18] ),
    .X(_04465_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(\u_rf.reg2_q[18] ),
    .A1(_04465_),
    .S(_04449_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _09408_ (.A(_04466_),
    .X(_00018_));
 sky130_fd_sc_hd__clkbuf_2 _09409_ (.A(\u_decod.rf_ff_res_data_i[19] ),
    .X(_04467_));
 sky130_fd_sc_hd__mux2_1 _09410_ (.A0(\u_rf.reg2_q[19] ),
    .A1(_04467_),
    .S(_04449_),
    .X(_04468_));
 sky130_fd_sc_hd__clkbuf_1 _09411_ (.A(_04468_),
    .X(_00019_));
 sky130_fd_sc_hd__buf_2 _09412_ (.A(\u_decod.rf_ff_res_data_i[20] ),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_8 _09413_ (.A(_04427_),
    .X(_04470_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(\u_rf.reg2_q[20] ),
    .A1(_04469_),
    .S(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _09415_ (.A(_04471_),
    .X(_00020_));
 sky130_fd_sc_hd__buf_2 _09416_ (.A(\u_decod.rf_ff_res_data_i[21] ),
    .X(_04472_));
 sky130_fd_sc_hd__mux2_1 _09417_ (.A0(\u_rf.reg2_q[21] ),
    .A1(_04472_),
    .S(_04470_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _09418_ (.A(_04473_),
    .X(_00021_));
 sky130_fd_sc_hd__buf_2 _09419_ (.A(\u_decod.rf_ff_res_data_i[22] ),
    .X(_04474_));
 sky130_fd_sc_hd__mux2_1 _09420_ (.A0(\u_rf.reg2_q[22] ),
    .A1(_04474_),
    .S(_04470_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _09421_ (.A(_04475_),
    .X(_00022_));
 sky130_fd_sc_hd__buf_2 _09422_ (.A(\u_decod.rf_ff_res_data_i[23] ),
    .X(_04476_));
 sky130_fd_sc_hd__mux2_1 _09423_ (.A0(\u_rf.reg2_q[23] ),
    .A1(_04476_),
    .S(_04470_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _09424_ (.A(_04477_),
    .X(_00023_));
 sky130_fd_sc_hd__buf_2 _09425_ (.A(\u_decod.rf_ff_res_data_i[24] ),
    .X(_04478_));
 sky130_fd_sc_hd__mux2_1 _09426_ (.A0(\u_rf.reg2_q[24] ),
    .A1(_04478_),
    .S(_04470_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _09427_ (.A(_04479_),
    .X(_00024_));
 sky130_fd_sc_hd__buf_2 _09428_ (.A(\u_decod.rf_ff_res_data_i[25] ),
    .X(_04480_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(\u_rf.reg2_q[25] ),
    .A1(_04480_),
    .S(_04470_),
    .X(_04481_));
 sky130_fd_sc_hd__clkbuf_1 _09430_ (.A(_04481_),
    .X(_00025_));
 sky130_fd_sc_hd__buf_2 _09431_ (.A(\u_decod.rf_ff_res_data_i[26] ),
    .X(_04482_));
 sky130_fd_sc_hd__mux2_1 _09432_ (.A0(\u_rf.reg2_q[26] ),
    .A1(_04482_),
    .S(_04470_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _09433_ (.A(_04483_),
    .X(_00026_));
 sky130_fd_sc_hd__buf_2 _09434_ (.A(\u_decod.rf_ff_res_data_i[27] ),
    .X(_04484_));
 sky130_fd_sc_hd__mux2_1 _09435_ (.A0(\u_rf.reg2_q[27] ),
    .A1(_04484_),
    .S(_04470_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _09436_ (.A(_04485_),
    .X(_00027_));
 sky130_fd_sc_hd__buf_2 _09437_ (.A(\u_decod.rf_ff_res_data_i[28] ),
    .X(_04486_));
 sky130_fd_sc_hd__mux2_1 _09438_ (.A0(\u_rf.reg2_q[28] ),
    .A1(_04486_),
    .S(_04470_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _09439_ (.A(_04487_),
    .X(_00028_));
 sky130_fd_sc_hd__buf_2 _09440_ (.A(\u_decod.rf_ff_res_data_i[29] ),
    .X(_04488_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(\u_rf.reg2_q[29] ),
    .A1(_04488_),
    .S(_04470_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _09442_ (.A(_04489_),
    .X(_00029_));
 sky130_fd_sc_hd__buf_2 _09443_ (.A(\u_decod.rf_ff_res_data_i[30] ),
    .X(_04490_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(\u_rf.reg2_q[30] ),
    .A1(_04490_),
    .S(_04427_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _09445_ (.A(_04491_),
    .X(_00030_));
 sky130_fd_sc_hd__buf_2 _09446_ (.A(\u_decod.rf_ff_res_data_i[31] ),
    .X(_04492_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(\u_rf.reg2_q[31] ),
    .A1(_04492_),
    .S(_04427_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _09448_ (.A(_04493_),
    .X(_00031_));
 sky130_fd_sc_hd__or4_2 _09449_ (.A(_01534_),
    .B(_04424_),
    .C(_01531_),
    .D(_01536_),
    .X(_04494_));
 sky130_fd_sc_hd__nor2_2 _09450_ (.A(_04423_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__clkbuf_8 _09451_ (.A(_04495_),
    .X(_04496_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(\u_rf.reg1_q[0] ),
    .A1(_04421_),
    .S(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _09453_ (.A(_04497_),
    .X(_00032_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(\u_rf.reg1_q[1] ),
    .A1(_04430_),
    .S(_04496_),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_1 _09455_ (.A(_04498_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _09456_ (.A0(\u_rf.reg1_q[2] ),
    .A1(_04432_),
    .S(_04496_),
    .X(_04499_));
 sky130_fd_sc_hd__clkbuf_1 _09457_ (.A(_04499_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(\u_rf.reg1_q[3] ),
    .A1(_04434_),
    .S(_04496_),
    .X(_04500_));
 sky130_fd_sc_hd__clkbuf_1 _09459_ (.A(_04500_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(\u_rf.reg1_q[4] ),
    .A1(_04436_),
    .S(_04496_),
    .X(_04501_));
 sky130_fd_sc_hd__clkbuf_1 _09461_ (.A(_04501_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(\u_rf.reg1_q[5] ),
    .A1(_04438_),
    .S(_04496_),
    .X(_04502_));
 sky130_fd_sc_hd__clkbuf_1 _09463_ (.A(_04502_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(\u_rf.reg1_q[6] ),
    .A1(_04440_),
    .S(_04496_),
    .X(_04503_));
 sky130_fd_sc_hd__clkbuf_1 _09465_ (.A(_04503_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(\u_rf.reg1_q[7] ),
    .A1(_04442_),
    .S(_04496_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _09467_ (.A(_04504_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _09468_ (.A0(\u_rf.reg1_q[8] ),
    .A1(_04444_),
    .S(_04496_),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_1 _09469_ (.A(_04505_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _09470_ (.A0(\u_rf.reg1_q[9] ),
    .A1(_04446_),
    .S(_04496_),
    .X(_04506_));
 sky130_fd_sc_hd__clkbuf_1 _09471_ (.A(_04506_),
    .X(_00041_));
 sky130_fd_sc_hd__buf_6 _09472_ (.A(_04495_),
    .X(_04507_));
 sky130_fd_sc_hd__mux2_1 _09473_ (.A0(\u_rf.reg1_q[10] ),
    .A1(_04448_),
    .S(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__clkbuf_1 _09474_ (.A(_04508_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(\u_rf.reg1_q[11] ),
    .A1(_04451_),
    .S(_04507_),
    .X(_04509_));
 sky130_fd_sc_hd__clkbuf_1 _09476_ (.A(_04509_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(\u_rf.reg1_q[12] ),
    .A1(_04453_),
    .S(_04507_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _09478_ (.A(_04510_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _09479_ (.A0(\u_rf.reg1_q[13] ),
    .A1(_04455_),
    .S(_04507_),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_1 _09480_ (.A(_04511_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(\u_rf.reg1_q[14] ),
    .A1(_04457_),
    .S(_04507_),
    .X(_04512_));
 sky130_fd_sc_hd__clkbuf_1 _09482_ (.A(_04512_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _09483_ (.A0(\u_rf.reg1_q[15] ),
    .A1(_04459_),
    .S(_04507_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _09484_ (.A(_04513_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(\u_rf.reg1_q[16] ),
    .A1(_04461_),
    .S(_04507_),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_1 _09486_ (.A(_04514_),
    .X(_00048_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(\u_rf.reg1_q[17] ),
    .A1(_04463_),
    .S(_04507_),
    .X(_04515_));
 sky130_fd_sc_hd__clkbuf_1 _09488_ (.A(_04515_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _09489_ (.A0(\u_rf.reg1_q[18] ),
    .A1(_04465_),
    .S(_04507_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _09490_ (.A(_04516_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(\u_rf.reg1_q[19] ),
    .A1(_04467_),
    .S(_04507_),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_1 _09492_ (.A(_04517_),
    .X(_00051_));
 sky130_fd_sc_hd__clkbuf_8 _09493_ (.A(_04495_),
    .X(_04518_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(\u_rf.reg1_q[20] ),
    .A1(_04469_),
    .S(_04518_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _09495_ (.A(_04519_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _09496_ (.A0(\u_rf.reg1_q[21] ),
    .A1(_04472_),
    .S(_04518_),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_1 _09497_ (.A(_04520_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _09498_ (.A0(\u_rf.reg1_q[22] ),
    .A1(_04474_),
    .S(_04518_),
    .X(_04521_));
 sky130_fd_sc_hd__clkbuf_1 _09499_ (.A(_04521_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _09500_ (.A0(\u_rf.reg1_q[23] ),
    .A1(_04476_),
    .S(_04518_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _09501_ (.A(_04522_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _09502_ (.A0(\u_rf.reg1_q[24] ),
    .A1(_04478_),
    .S(_04518_),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_1 _09503_ (.A(_04523_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _09504_ (.A0(\u_rf.reg1_q[25] ),
    .A1(_04480_),
    .S(_04518_),
    .X(_04524_));
 sky130_fd_sc_hd__clkbuf_1 _09505_ (.A(_04524_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(\u_rf.reg1_q[26] ),
    .A1(_04482_),
    .S(_04518_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_1 _09507_ (.A(_04525_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _09508_ (.A0(\u_rf.reg1_q[27] ),
    .A1(_04484_),
    .S(_04518_),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_1 _09509_ (.A(_04526_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _09510_ (.A0(\u_rf.reg1_q[28] ),
    .A1(_04486_),
    .S(_04518_),
    .X(_04527_));
 sky130_fd_sc_hd__clkbuf_1 _09511_ (.A(_04527_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _09512_ (.A0(\u_rf.reg1_q[29] ),
    .A1(_04488_),
    .S(_04518_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _09513_ (.A(_04528_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _09514_ (.A0(\u_rf.reg1_q[30] ),
    .A1(_04490_),
    .S(_04495_),
    .X(_04529_));
 sky130_fd_sc_hd__clkbuf_1 _09515_ (.A(_04529_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _09516_ (.A0(\u_rf.reg1_q[31] ),
    .A1(_04492_),
    .S(_04495_),
    .X(_04530_));
 sky130_fd_sc_hd__clkbuf_1 _09517_ (.A(_04530_),
    .X(_00063_));
 sky130_fd_sc_hd__or4_2 _09518_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_04424_),
    .C(_01531_),
    .D(_01536_),
    .X(_04531_));
 sky130_fd_sc_hd__nor2_2 _09519_ (.A(_04423_),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__clkbuf_8 _09520_ (.A(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(\u_rf.reg0_q[0] ),
    .A1(_04421_),
    .S(_04533_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _09522_ (.A(_04534_),
    .X(_00064_));
 sky130_fd_sc_hd__mux2_1 _09523_ (.A0(\u_rf.reg0_q[1] ),
    .A1(_04430_),
    .S(_04533_),
    .X(_04535_));
 sky130_fd_sc_hd__clkbuf_1 _09524_ (.A(_04535_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(\u_rf.reg0_q[2] ),
    .A1(_04432_),
    .S(_04533_),
    .X(_04536_));
 sky130_fd_sc_hd__clkbuf_1 _09526_ (.A(_04536_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _09527_ (.A0(\u_rf.reg0_q[3] ),
    .A1(_04434_),
    .S(_04533_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _09528_ (.A(_04537_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(\u_rf.reg0_q[4] ),
    .A1(_04436_),
    .S(_04533_),
    .X(_04538_));
 sky130_fd_sc_hd__clkbuf_1 _09530_ (.A(_04538_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(\u_rf.reg0_q[5] ),
    .A1(_04438_),
    .S(_04533_),
    .X(_04539_));
 sky130_fd_sc_hd__clkbuf_1 _09532_ (.A(_04539_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _09533_ (.A0(\u_rf.reg0_q[6] ),
    .A1(_04440_),
    .S(_04533_),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_1 _09534_ (.A(_04540_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(\u_rf.reg0_q[7] ),
    .A1(_04442_),
    .S(_04533_),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_1 _09536_ (.A(_04541_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(\u_rf.reg0_q[8] ),
    .A1(_04444_),
    .S(_04533_),
    .X(_04542_));
 sky130_fd_sc_hd__clkbuf_1 _09538_ (.A(_04542_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _09539_ (.A0(\u_rf.reg0_q[9] ),
    .A1(_04446_),
    .S(_04533_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _09540_ (.A(_04543_),
    .X(_00073_));
 sky130_fd_sc_hd__buf_6 _09541_ (.A(_04532_),
    .X(_04544_));
 sky130_fd_sc_hd__mux2_1 _09542_ (.A0(\u_rf.reg0_q[10] ),
    .A1(_04448_),
    .S(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__clkbuf_1 _09543_ (.A(_04545_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _09544_ (.A0(\u_rf.reg0_q[11] ),
    .A1(_04451_),
    .S(_04544_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _09545_ (.A(_04546_),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _09546_ (.A0(\u_rf.reg0_q[12] ),
    .A1(_04453_),
    .S(_04544_),
    .X(_04547_));
 sky130_fd_sc_hd__clkbuf_1 _09547_ (.A(_04547_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _09548_ (.A0(\u_rf.reg0_q[13] ),
    .A1(_04455_),
    .S(_04544_),
    .X(_04548_));
 sky130_fd_sc_hd__clkbuf_1 _09549_ (.A(_04548_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _09550_ (.A0(\u_rf.reg0_q[14] ),
    .A1(_04457_),
    .S(_04544_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _09551_ (.A(_04549_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _09552_ (.A0(\u_rf.reg0_q[15] ),
    .A1(_04459_),
    .S(_04544_),
    .X(_04550_));
 sky130_fd_sc_hd__clkbuf_1 _09553_ (.A(_04550_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _09554_ (.A0(\u_rf.reg0_q[16] ),
    .A1(_04461_),
    .S(_04544_),
    .X(_04551_));
 sky130_fd_sc_hd__clkbuf_1 _09555_ (.A(_04551_),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _09556_ (.A0(\u_rf.reg0_q[17] ),
    .A1(_04463_),
    .S(_04544_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _09557_ (.A(_04552_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _09558_ (.A0(\u_rf.reg0_q[18] ),
    .A1(_04465_),
    .S(_04544_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_1 _09559_ (.A(_04553_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _09560_ (.A0(\u_rf.reg0_q[19] ),
    .A1(_04467_),
    .S(_04544_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _09561_ (.A(_04554_),
    .X(_00083_));
 sky130_fd_sc_hd__clkbuf_8 _09562_ (.A(_04532_),
    .X(_04555_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(\u_rf.reg0_q[20] ),
    .A1(_04469_),
    .S(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _09564_ (.A(_04556_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(\u_rf.reg0_q[21] ),
    .A1(_04472_),
    .S(_04555_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _09566_ (.A(_04557_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(\u_rf.reg0_q[22] ),
    .A1(_04474_),
    .S(_04555_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _09568_ (.A(_04558_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(\u_rf.reg0_q[23] ),
    .A1(_04476_),
    .S(_04555_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _09570_ (.A(_04559_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(\u_rf.reg0_q[24] ),
    .A1(_04478_),
    .S(_04555_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _09572_ (.A(_04560_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(\u_rf.reg0_q[25] ),
    .A1(_04480_),
    .S(_04555_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _09574_ (.A(_04561_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(\u_rf.reg0_q[26] ),
    .A1(_04482_),
    .S(_04555_),
    .X(_04562_));
 sky130_fd_sc_hd__clkbuf_1 _09576_ (.A(_04562_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _09577_ (.A0(\u_rf.reg0_q[27] ),
    .A1(_04484_),
    .S(_04555_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _09578_ (.A(_04563_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(\u_rf.reg0_q[28] ),
    .A1(_04486_),
    .S(_04555_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _09580_ (.A(_04564_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(\u_rf.reg0_q[29] ),
    .A1(_04488_),
    .S(_04555_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _09582_ (.A(_04565_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(\u_rf.reg0_q[30] ),
    .A1(_04490_),
    .S(_04532_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _09584_ (.A(_04566_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(\u_rf.reg0_q[31] ),
    .A1(_04492_),
    .S(_04532_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _09586_ (.A(_04567_),
    .X(_00095_));
 sky130_fd_sc_hd__nand2_2 _09587_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_04424_),
    .Y(_04568_));
 sky130_fd_sc_hd__or3_2 _09588_ (.A(_01531_),
    .B(_01536_),
    .C(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__nor2_4 _09589_ (.A(_04423_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__clkbuf_8 _09590_ (.A(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _09591_ (.A0(\u_rf.reg3_q[0] ),
    .A1(_04421_),
    .S(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _09592_ (.A(_04572_),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(\u_rf.reg3_q[1] ),
    .A1(_04430_),
    .S(_04571_),
    .X(_04573_));
 sky130_fd_sc_hd__clkbuf_1 _09594_ (.A(_04573_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _09595_ (.A0(\u_rf.reg3_q[2] ),
    .A1(_04432_),
    .S(_04571_),
    .X(_04574_));
 sky130_fd_sc_hd__clkbuf_1 _09596_ (.A(_04574_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(\u_rf.reg3_q[3] ),
    .A1(_04434_),
    .S(_04571_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_1 _09598_ (.A(_04575_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(\u_rf.reg3_q[4] ),
    .A1(_04436_),
    .S(_04571_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _09600_ (.A(_04576_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(\u_rf.reg3_q[5] ),
    .A1(_04438_),
    .S(_04571_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _09602_ (.A(_04577_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _09603_ (.A0(\u_rf.reg3_q[6] ),
    .A1(_04440_),
    .S(_04571_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _09604_ (.A(_04578_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(\u_rf.reg3_q[7] ),
    .A1(_04442_),
    .S(_04571_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _09606_ (.A(_04579_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _09607_ (.A0(\u_rf.reg3_q[8] ),
    .A1(_04444_),
    .S(_04571_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _09608_ (.A(_04580_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(\u_rf.reg3_q[9] ),
    .A1(_04446_),
    .S(_04571_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_1 _09610_ (.A(_04581_),
    .X(_00105_));
 sky130_fd_sc_hd__buf_6 _09611_ (.A(_04570_),
    .X(_04582_));
 sky130_fd_sc_hd__mux2_1 _09612_ (.A0(\u_rf.reg3_q[10] ),
    .A1(_04448_),
    .S(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _09613_ (.A(_04583_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _09614_ (.A0(\u_rf.reg3_q[11] ),
    .A1(_04451_),
    .S(_04582_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_1 _09615_ (.A(_04584_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _09616_ (.A0(\u_rf.reg3_q[12] ),
    .A1(_04453_),
    .S(_04582_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _09617_ (.A(_04585_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _09618_ (.A0(\u_rf.reg3_q[13] ),
    .A1(_04455_),
    .S(_04582_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _09619_ (.A(_04586_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _09620_ (.A0(\u_rf.reg3_q[14] ),
    .A1(_04457_),
    .S(_04582_),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_1 _09621_ (.A(_04587_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _09622_ (.A0(\u_rf.reg3_q[15] ),
    .A1(_04459_),
    .S(_04582_),
    .X(_04588_));
 sky130_fd_sc_hd__clkbuf_1 _09623_ (.A(_04588_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(\u_rf.reg3_q[16] ),
    .A1(_04461_),
    .S(_04582_),
    .X(_04589_));
 sky130_fd_sc_hd__clkbuf_1 _09625_ (.A(_04589_),
    .X(_00112_));
 sky130_fd_sc_hd__mux2_1 _09626_ (.A0(\u_rf.reg3_q[17] ),
    .A1(_04463_),
    .S(_04582_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _09627_ (.A(_04590_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _09628_ (.A0(\u_rf.reg3_q[18] ),
    .A1(_04465_),
    .S(_04582_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _09629_ (.A(_04591_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(\u_rf.reg3_q[19] ),
    .A1(_04467_),
    .S(_04582_),
    .X(_04592_));
 sky130_fd_sc_hd__clkbuf_1 _09631_ (.A(_04592_),
    .X(_00115_));
 sky130_fd_sc_hd__clkbuf_8 _09632_ (.A(_04570_),
    .X(_04593_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(\u_rf.reg3_q[20] ),
    .A1(_04469_),
    .S(_04593_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _09634_ (.A(_04594_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(\u_rf.reg3_q[21] ),
    .A1(_04472_),
    .S(_04593_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _09636_ (.A(_04595_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(\u_rf.reg3_q[22] ),
    .A1(_04474_),
    .S(_04593_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _09638_ (.A(_04596_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(\u_rf.reg3_q[23] ),
    .A1(_04476_),
    .S(_04593_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _09640_ (.A(_04597_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(\u_rf.reg3_q[24] ),
    .A1(_04478_),
    .S(_04593_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _09642_ (.A(_04598_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _09643_ (.A0(\u_rf.reg3_q[25] ),
    .A1(_04480_),
    .S(_04593_),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_1 _09644_ (.A(_04599_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(\u_rf.reg3_q[26] ),
    .A1(_04482_),
    .S(_04593_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _09646_ (.A(_04600_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(\u_rf.reg3_q[27] ),
    .A1(_04484_),
    .S(_04593_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _09648_ (.A(_04601_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(\u_rf.reg3_q[28] ),
    .A1(_04486_),
    .S(_04593_),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_1 _09650_ (.A(_04602_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(\u_rf.reg3_q[29] ),
    .A1(_04488_),
    .S(_04593_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_04603_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(\u_rf.reg3_q[30] ),
    .A1(_04490_),
    .S(_04570_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _09654_ (.A(_04604_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(\u_rf.reg3_q[31] ),
    .A1(_04492_),
    .S(_04570_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _09656_ (.A(_04605_),
    .X(_00127_));
 sky130_fd_sc_hd__or4_2 _09657_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_04424_),
    .C(_01532_),
    .D(_01536_),
    .X(_04606_));
 sky130_fd_sc_hd__nor2_4 _09658_ (.A(_04423_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__buf_6 _09659_ (.A(_04607_),
    .X(_04608_));
 sky130_fd_sc_hd__mux2_1 _09660_ (.A0(\u_rf.reg4_q[0] ),
    .A1(_04421_),
    .S(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__clkbuf_1 _09661_ (.A(_04609_),
    .X(_00128_));
 sky130_fd_sc_hd__mux2_1 _09662_ (.A0(\u_rf.reg4_q[1] ),
    .A1(_04430_),
    .S(_04608_),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_1 _09663_ (.A(_04610_),
    .X(_00129_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(\u_rf.reg4_q[2] ),
    .A1(_04432_),
    .S(_04608_),
    .X(_04611_));
 sky130_fd_sc_hd__clkbuf_1 _09665_ (.A(_04611_),
    .X(_00130_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(\u_rf.reg4_q[3] ),
    .A1(_04434_),
    .S(_04608_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _09667_ (.A(_04612_),
    .X(_00131_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(\u_rf.reg4_q[4] ),
    .A1(_04436_),
    .S(_04608_),
    .X(_04613_));
 sky130_fd_sc_hd__clkbuf_1 _09669_ (.A(_04613_),
    .X(_00132_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(\u_rf.reg4_q[5] ),
    .A1(_04438_),
    .S(_04608_),
    .X(_04614_));
 sky130_fd_sc_hd__clkbuf_1 _09671_ (.A(_04614_),
    .X(_00133_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(\u_rf.reg4_q[6] ),
    .A1(_04440_),
    .S(_04608_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _09673_ (.A(_04615_),
    .X(_00134_));
 sky130_fd_sc_hd__mux2_1 _09674_ (.A0(\u_rf.reg4_q[7] ),
    .A1(_04442_),
    .S(_04608_),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_1 _09675_ (.A(_04616_),
    .X(_00135_));
 sky130_fd_sc_hd__mux2_1 _09676_ (.A0(\u_rf.reg4_q[8] ),
    .A1(_04444_),
    .S(_04608_),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_1 _09677_ (.A(_04617_),
    .X(_00136_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(\u_rf.reg4_q[9] ),
    .A1(_04446_),
    .S(_04608_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_1 _09679_ (.A(_04618_),
    .X(_00137_));
 sky130_fd_sc_hd__buf_6 _09680_ (.A(_04607_),
    .X(_04619_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(\u_rf.reg4_q[10] ),
    .A1(_04448_),
    .S(_04619_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _09682_ (.A(_04620_),
    .X(_00138_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(\u_rf.reg4_q[11] ),
    .A1(_04451_),
    .S(_04619_),
    .X(_04621_));
 sky130_fd_sc_hd__clkbuf_1 _09684_ (.A(_04621_),
    .X(_00139_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(\u_rf.reg4_q[12] ),
    .A1(_04453_),
    .S(_04619_),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_1 _09686_ (.A(_04622_),
    .X(_00140_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(\u_rf.reg4_q[13] ),
    .A1(_04455_),
    .S(_04619_),
    .X(_04623_));
 sky130_fd_sc_hd__clkbuf_1 _09688_ (.A(_04623_),
    .X(_00141_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(\u_rf.reg4_q[14] ),
    .A1(_04457_),
    .S(_04619_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _09690_ (.A(_04624_),
    .X(_00142_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(\u_rf.reg4_q[15] ),
    .A1(_04459_),
    .S(_04619_),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _09692_ (.A(_04625_),
    .X(_00143_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(\u_rf.reg4_q[16] ),
    .A1(_04461_),
    .S(_04619_),
    .X(_04626_));
 sky130_fd_sc_hd__clkbuf_1 _09694_ (.A(_04626_),
    .X(_00144_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(\u_rf.reg4_q[17] ),
    .A1(_04463_),
    .S(_04619_),
    .X(_04627_));
 sky130_fd_sc_hd__clkbuf_1 _09696_ (.A(_04627_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _09697_ (.A0(\u_rf.reg4_q[18] ),
    .A1(_04465_),
    .S(_04619_),
    .X(_04628_));
 sky130_fd_sc_hd__clkbuf_1 _09698_ (.A(_04628_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(\u_rf.reg4_q[19] ),
    .A1(_04467_),
    .S(_04619_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _09700_ (.A(_04629_),
    .X(_00147_));
 sky130_fd_sc_hd__clkbuf_8 _09701_ (.A(_04607_),
    .X(_04630_));
 sky130_fd_sc_hd__mux2_1 _09702_ (.A0(\u_rf.reg4_q[20] ),
    .A1(_04469_),
    .S(_04630_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _09703_ (.A(_04631_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _09704_ (.A0(\u_rf.reg4_q[21] ),
    .A1(_04472_),
    .S(_04630_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _09705_ (.A(_04632_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _09706_ (.A0(\u_rf.reg4_q[22] ),
    .A1(_04474_),
    .S(_04630_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _09707_ (.A(_04633_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _09708_ (.A0(\u_rf.reg4_q[23] ),
    .A1(_04476_),
    .S(_04630_),
    .X(_04634_));
 sky130_fd_sc_hd__clkbuf_1 _09709_ (.A(_04634_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _09710_ (.A0(\u_rf.reg4_q[24] ),
    .A1(_04478_),
    .S(_04630_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _09711_ (.A(_04635_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(\u_rf.reg4_q[25] ),
    .A1(_04480_),
    .S(_04630_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _09713_ (.A(_04636_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _09714_ (.A0(\u_rf.reg4_q[26] ),
    .A1(_04482_),
    .S(_04630_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _09715_ (.A(_04637_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _09716_ (.A0(\u_rf.reg4_q[27] ),
    .A1(_04484_),
    .S(_04630_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _09717_ (.A(_04638_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(\u_rf.reg4_q[28] ),
    .A1(_04486_),
    .S(_04630_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _09719_ (.A(_04639_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(\u_rf.reg4_q[29] ),
    .A1(_04488_),
    .S(_04630_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_1 _09721_ (.A(_04640_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(\u_rf.reg4_q[30] ),
    .A1(_04490_),
    .S(_04607_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _09723_ (.A(_04641_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(\u_rf.reg4_q[31] ),
    .A1(_04492_),
    .S(_04607_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _09725_ (.A(_04642_),
    .X(_00159_));
 sky130_fd_sc_hd__and2_1 _09726_ (.A(_01539_),
    .B(\u_decod.rf_write_v_q_i ),
    .X(_04643_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(_01534_),
    .B(_04424_),
    .Y(_04644_));
 sky130_fd_sc_hd__nor2_1 _09728_ (.A(_01532_),
    .B(_01536_),
    .Y(_04645_));
 sky130_fd_sc_hd__and3_4 _09729_ (.A(_04643_),
    .B(_04644_),
    .C(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__clkbuf_8 _09730_ (.A(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__mux2_1 _09731_ (.A0(\u_rf.reg5_q[0] ),
    .A1(_04421_),
    .S(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__clkbuf_1 _09732_ (.A(_04648_),
    .X(_00160_));
 sky130_fd_sc_hd__mux2_1 _09733_ (.A0(\u_rf.reg5_q[1] ),
    .A1(_04430_),
    .S(_04647_),
    .X(_04649_));
 sky130_fd_sc_hd__clkbuf_1 _09734_ (.A(_04649_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _09735_ (.A0(\u_rf.reg5_q[2] ),
    .A1(_04432_),
    .S(_04647_),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _09736_ (.A(_04650_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(\u_rf.reg5_q[3] ),
    .A1(_04434_),
    .S(_04647_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_1 _09738_ (.A(_04651_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _09739_ (.A0(\u_rf.reg5_q[4] ),
    .A1(_04436_),
    .S(_04647_),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_1 _09740_ (.A(_04652_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _09741_ (.A0(\u_rf.reg5_q[5] ),
    .A1(_04438_),
    .S(_04647_),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_1 _09742_ (.A(_04653_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(\u_rf.reg5_q[6] ),
    .A1(_04440_),
    .S(_04647_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_04654_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _09745_ (.A0(\u_rf.reg5_q[7] ),
    .A1(_04442_),
    .S(_04647_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_1 _09746_ (.A(_04655_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _09747_ (.A0(\u_rf.reg5_q[8] ),
    .A1(_04444_),
    .S(_04647_),
    .X(_04656_));
 sky130_fd_sc_hd__clkbuf_1 _09748_ (.A(_04656_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(\u_rf.reg5_q[9] ),
    .A1(_04446_),
    .S(_04647_),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(_04657_),
    .X(_00169_));
 sky130_fd_sc_hd__buf_6 _09751_ (.A(_04646_),
    .X(_04658_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(\u_rf.reg5_q[10] ),
    .A1(_04448_),
    .S(_04658_),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_1 _09753_ (.A(_04659_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _09754_ (.A0(\u_rf.reg5_q[11] ),
    .A1(_04451_),
    .S(_04658_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _09755_ (.A(_04660_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _09756_ (.A0(\u_rf.reg5_q[12] ),
    .A1(_04453_),
    .S(_04658_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _09757_ (.A(_04661_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(\u_rf.reg5_q[13] ),
    .A1(_04455_),
    .S(_04658_),
    .X(_04662_));
 sky130_fd_sc_hd__clkbuf_1 _09759_ (.A(_04662_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _09760_ (.A0(\u_rf.reg5_q[14] ),
    .A1(_04457_),
    .S(_04658_),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _09761_ (.A(_04663_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _09762_ (.A0(\u_rf.reg5_q[15] ),
    .A1(_04459_),
    .S(_04658_),
    .X(_04664_));
 sky130_fd_sc_hd__clkbuf_1 _09763_ (.A(_04664_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(\u_rf.reg5_q[16] ),
    .A1(_04461_),
    .S(_04658_),
    .X(_04665_));
 sky130_fd_sc_hd__clkbuf_1 _09765_ (.A(_04665_),
    .X(_00176_));
 sky130_fd_sc_hd__mux2_1 _09766_ (.A0(\u_rf.reg5_q[17] ),
    .A1(_04463_),
    .S(_04658_),
    .X(_04666_));
 sky130_fd_sc_hd__clkbuf_1 _09767_ (.A(_04666_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _09768_ (.A0(\u_rf.reg5_q[18] ),
    .A1(_04465_),
    .S(_04658_),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _09769_ (.A(_04667_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(\u_rf.reg5_q[19] ),
    .A1(_04467_),
    .S(_04658_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_1 _09771_ (.A(_04668_),
    .X(_00179_));
 sky130_fd_sc_hd__buf_6 _09772_ (.A(_04646_),
    .X(_04669_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(\u_rf.reg5_q[20] ),
    .A1(_04469_),
    .S(_04669_),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_1 _09774_ (.A(_04670_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _09775_ (.A0(\u_rf.reg5_q[21] ),
    .A1(_04472_),
    .S(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _09776_ (.A(_04671_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _09777_ (.A0(\u_rf.reg5_q[22] ),
    .A1(_04474_),
    .S(_04669_),
    .X(_04672_));
 sky130_fd_sc_hd__clkbuf_1 _09778_ (.A(_04672_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(\u_rf.reg5_q[23] ),
    .A1(_04476_),
    .S(_04669_),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _09780_ (.A(_04673_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _09781_ (.A0(\u_rf.reg5_q[24] ),
    .A1(_04478_),
    .S(_04669_),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_1 _09782_ (.A(_04674_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _09783_ (.A0(\u_rf.reg5_q[25] ),
    .A1(_04480_),
    .S(_04669_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _09784_ (.A(_04675_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(\u_rf.reg5_q[26] ),
    .A1(_04482_),
    .S(_04669_),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_04676_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(\u_rf.reg5_q[27] ),
    .A1(_04484_),
    .S(_04669_),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_04677_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(\u_rf.reg5_q[28] ),
    .A1(_04486_),
    .S(_04669_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _09790_ (.A(_04678_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(\u_rf.reg5_q[29] ),
    .A1(_04488_),
    .S(_04669_),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _09792_ (.A(_04679_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(\u_rf.reg5_q[30] ),
    .A1(_04490_),
    .S(_04646_),
    .X(_04680_));
 sky130_fd_sc_hd__clkbuf_1 _09794_ (.A(_04680_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(\u_rf.reg5_q[31] ),
    .A1(_04492_),
    .S(_04646_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _09796_ (.A(_04681_),
    .X(_00191_));
 sky130_fd_sc_hd__nor2_1 _09797_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_01542_),
    .Y(_04682_));
 sky130_fd_sc_hd__and3_4 _09798_ (.A(_04643_),
    .B(_04682_),
    .C(_04645_),
    .X(_04683_));
 sky130_fd_sc_hd__buf_6 _09799_ (.A(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__mux2_1 _09800_ (.A0(\u_rf.reg6_q[0] ),
    .A1(_04421_),
    .S(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__clkbuf_1 _09801_ (.A(_04685_),
    .X(_00192_));
 sky130_fd_sc_hd__mux2_1 _09802_ (.A0(\u_rf.reg6_q[1] ),
    .A1(_04430_),
    .S(_04684_),
    .X(_04686_));
 sky130_fd_sc_hd__clkbuf_1 _09803_ (.A(_04686_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _09804_ (.A0(\u_rf.reg6_q[2] ),
    .A1(_04432_),
    .S(_04684_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _09805_ (.A(_04687_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _09806_ (.A0(\u_rf.reg6_q[3] ),
    .A1(_04434_),
    .S(_04684_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _09807_ (.A(_04688_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _09808_ (.A0(\u_rf.reg6_q[4] ),
    .A1(_04436_),
    .S(_04684_),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_1 _09809_ (.A(_04689_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _09810_ (.A0(\u_rf.reg6_q[5] ),
    .A1(_04438_),
    .S(_04684_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _09811_ (.A(_04690_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _09812_ (.A0(\u_rf.reg6_q[6] ),
    .A1(_04440_),
    .S(_04684_),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_1 _09813_ (.A(_04691_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _09814_ (.A0(\u_rf.reg6_q[7] ),
    .A1(_04442_),
    .S(_04684_),
    .X(_04692_));
 sky130_fd_sc_hd__clkbuf_1 _09815_ (.A(_04692_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _09816_ (.A0(\u_rf.reg6_q[8] ),
    .A1(_04444_),
    .S(_04684_),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _09817_ (.A(_04693_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _09818_ (.A0(\u_rf.reg6_q[9] ),
    .A1(_04446_),
    .S(_04684_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _09819_ (.A(_04694_),
    .X(_00201_));
 sky130_fd_sc_hd__clkbuf_8 _09820_ (.A(_04683_),
    .X(_04695_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(\u_rf.reg6_q[10] ),
    .A1(_04448_),
    .S(_04695_),
    .X(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _09822_ (.A(_04696_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(\u_rf.reg6_q[11] ),
    .A1(_04451_),
    .S(_04695_),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_1 _09824_ (.A(_04697_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(\u_rf.reg6_q[12] ),
    .A1(_04453_),
    .S(_04695_),
    .X(_04698_));
 sky130_fd_sc_hd__clkbuf_1 _09826_ (.A(_04698_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(\u_rf.reg6_q[13] ),
    .A1(_04455_),
    .S(_04695_),
    .X(_04699_));
 sky130_fd_sc_hd__clkbuf_1 _09828_ (.A(_04699_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _09829_ (.A0(\u_rf.reg6_q[14] ),
    .A1(_04457_),
    .S(_04695_),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_1 _09830_ (.A(_04700_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(\u_rf.reg6_q[15] ),
    .A1(_04459_),
    .S(_04695_),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _09832_ (.A(_04701_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(\u_rf.reg6_q[16] ),
    .A1(_04461_),
    .S(_04695_),
    .X(_04702_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_04702_),
    .X(_00208_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(\u_rf.reg6_q[17] ),
    .A1(_04463_),
    .S(_04695_),
    .X(_04703_));
 sky130_fd_sc_hd__clkbuf_1 _09836_ (.A(_04703_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(\u_rf.reg6_q[18] ),
    .A1(_04465_),
    .S(_04695_),
    .X(_04704_));
 sky130_fd_sc_hd__clkbuf_1 _09838_ (.A(_04704_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _09839_ (.A0(\u_rf.reg6_q[19] ),
    .A1(_04467_),
    .S(_04695_),
    .X(_04705_));
 sky130_fd_sc_hd__clkbuf_1 _09840_ (.A(_04705_),
    .X(_00211_));
 sky130_fd_sc_hd__clkbuf_8 _09841_ (.A(_04683_),
    .X(_04706_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(\u_rf.reg6_q[20] ),
    .A1(_04469_),
    .S(_04706_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _09843_ (.A(_04707_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(\u_rf.reg6_q[21] ),
    .A1(_04472_),
    .S(_04706_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _09845_ (.A(_04708_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _09846_ (.A0(\u_rf.reg6_q[22] ),
    .A1(_04474_),
    .S(_04706_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _09847_ (.A(_04709_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(\u_rf.reg6_q[23] ),
    .A1(_04476_),
    .S(_04706_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _09849_ (.A(_04710_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(\u_rf.reg6_q[24] ),
    .A1(_04478_),
    .S(_04706_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _09851_ (.A(_04711_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(\u_rf.reg6_q[25] ),
    .A1(_04480_),
    .S(_04706_),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_1 _09853_ (.A(_04712_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _09854_ (.A0(\u_rf.reg6_q[26] ),
    .A1(_04482_),
    .S(_04706_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _09855_ (.A(_04713_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _09856_ (.A0(\u_rf.reg6_q[27] ),
    .A1(_04484_),
    .S(_04706_),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _09857_ (.A(_04714_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(\u_rf.reg6_q[28] ),
    .A1(_04486_),
    .S(_04706_),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_1 _09859_ (.A(_04715_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(\u_rf.reg6_q[29] ),
    .A1(_04488_),
    .S(_04706_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_1 _09861_ (.A(_04716_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(\u_rf.reg6_q[30] ),
    .A1(_04490_),
    .S(_04683_),
    .X(_04717_));
 sky130_fd_sc_hd__clkbuf_1 _09863_ (.A(_04717_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _09864_ (.A0(\u_rf.reg6_q[31] ),
    .A1(_04492_),
    .S(_04683_),
    .X(_04718_));
 sky130_fd_sc_hd__clkbuf_1 _09865_ (.A(_04718_),
    .X(_00223_));
 sky130_fd_sc_hd__buf_2 _09866_ (.A(\u_decod.rf_ff_res_data_i[0] ),
    .X(_04719_));
 sky130_fd_sc_hd__or3b_1 _09867_ (.A(_04422_),
    .B(_04568_),
    .C_N(_04645_),
    .X(_04720_));
 sky130_fd_sc_hd__clkbuf_4 _09868_ (.A(_04720_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_8 _09869_ (.A(_04721_),
    .X(_04722_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(_04719_),
    .A1(\u_rf.reg7_q[0] ),
    .S(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__clkbuf_1 _09871_ (.A(_04723_),
    .X(_00224_));
 sky130_fd_sc_hd__buf_2 _09872_ (.A(\u_decod.rf_ff_res_data_i[1] ),
    .X(_04724_));
 sky130_fd_sc_hd__mux2_1 _09873_ (.A0(_04724_),
    .A1(\u_rf.reg7_q[1] ),
    .S(_04722_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _09874_ (.A(_04725_),
    .X(_00225_));
 sky130_fd_sc_hd__clkbuf_2 _09875_ (.A(\u_decod.rf_ff_res_data_i[2] ),
    .X(_04726_));
 sky130_fd_sc_hd__mux2_1 _09876_ (.A0(_04726_),
    .A1(\u_rf.reg7_q[2] ),
    .S(_04722_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _09877_ (.A(_04727_),
    .X(_00226_));
 sky130_fd_sc_hd__buf_2 _09878_ (.A(\u_decod.rf_ff_res_data_i[3] ),
    .X(_04728_));
 sky130_fd_sc_hd__mux2_1 _09879_ (.A0(_04728_),
    .A1(\u_rf.reg7_q[3] ),
    .S(_04722_),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_1 _09880_ (.A(_04729_),
    .X(_00227_));
 sky130_fd_sc_hd__clkbuf_2 _09881_ (.A(\u_decod.rf_ff_res_data_i[4] ),
    .X(_04730_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(_04730_),
    .A1(\u_rf.reg7_q[4] ),
    .S(_04722_),
    .X(_04731_));
 sky130_fd_sc_hd__clkbuf_1 _09883_ (.A(_04731_),
    .X(_00228_));
 sky130_fd_sc_hd__clkbuf_2 _09884_ (.A(\u_decod.rf_ff_res_data_i[5] ),
    .X(_04732_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(_04732_),
    .A1(\u_rf.reg7_q[5] ),
    .S(_04722_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _09886_ (.A(_04733_),
    .X(_00229_));
 sky130_fd_sc_hd__clkbuf_2 _09887_ (.A(\u_decod.rf_ff_res_data_i[6] ),
    .X(_04734_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(_04734_),
    .A1(\u_rf.reg7_q[6] ),
    .S(_04722_),
    .X(_04735_));
 sky130_fd_sc_hd__clkbuf_1 _09889_ (.A(_04735_),
    .X(_00230_));
 sky130_fd_sc_hd__clkbuf_2 _09890_ (.A(\u_decod.rf_ff_res_data_i[7] ),
    .X(_04736_));
 sky130_fd_sc_hd__mux2_1 _09891_ (.A0(_04736_),
    .A1(\u_rf.reg7_q[7] ),
    .S(_04722_),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_1 _09892_ (.A(_04737_),
    .X(_00231_));
 sky130_fd_sc_hd__clkbuf_2 _09893_ (.A(\u_decod.rf_ff_res_data_i[8] ),
    .X(_04738_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(_04738_),
    .A1(\u_rf.reg7_q[8] ),
    .S(_04722_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_1 _09895_ (.A(_04739_),
    .X(_00232_));
 sky130_fd_sc_hd__buf_2 _09896_ (.A(\u_decod.rf_ff_res_data_i[9] ),
    .X(_04740_));
 sky130_fd_sc_hd__mux2_1 _09897_ (.A0(_04740_),
    .A1(\u_rf.reg7_q[9] ),
    .S(_04722_),
    .X(_04741_));
 sky130_fd_sc_hd__clkbuf_1 _09898_ (.A(_04741_),
    .X(_00233_));
 sky130_fd_sc_hd__clkbuf_2 _09899_ (.A(\u_decod.rf_ff_res_data_i[10] ),
    .X(_04742_));
 sky130_fd_sc_hd__clkbuf_8 _09900_ (.A(_04721_),
    .X(_04743_));
 sky130_fd_sc_hd__mux2_1 _09901_ (.A0(_04742_),
    .A1(\u_rf.reg7_q[10] ),
    .S(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_1 _09902_ (.A(_04744_),
    .X(_00234_));
 sky130_fd_sc_hd__clkbuf_2 _09903_ (.A(\u_decod.rf_ff_res_data_i[11] ),
    .X(_04745_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(_04745_),
    .A1(\u_rf.reg7_q[11] ),
    .S(_04743_),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_1 _09905_ (.A(_04746_),
    .X(_00235_));
 sky130_fd_sc_hd__clkbuf_2 _09906_ (.A(\u_decod.rf_ff_res_data_i[12] ),
    .X(_04747_));
 sky130_fd_sc_hd__mux2_1 _09907_ (.A0(_04747_),
    .A1(\u_rf.reg7_q[12] ),
    .S(_04743_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _09908_ (.A(_04748_),
    .X(_00236_));
 sky130_fd_sc_hd__clkbuf_2 _09909_ (.A(\u_decod.rf_ff_res_data_i[13] ),
    .X(_04749_));
 sky130_fd_sc_hd__mux2_1 _09910_ (.A0(_04749_),
    .A1(\u_rf.reg7_q[13] ),
    .S(_04743_),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_1 _09911_ (.A(_04750_),
    .X(_00237_));
 sky130_fd_sc_hd__clkbuf_2 _09912_ (.A(\u_decod.rf_ff_res_data_i[14] ),
    .X(_04751_));
 sky130_fd_sc_hd__mux2_1 _09913_ (.A0(_04751_),
    .A1(\u_rf.reg7_q[14] ),
    .S(_04743_),
    .X(_04752_));
 sky130_fd_sc_hd__clkbuf_1 _09914_ (.A(_04752_),
    .X(_00238_));
 sky130_fd_sc_hd__clkbuf_2 _09915_ (.A(\u_decod.rf_ff_res_data_i[15] ),
    .X(_04753_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(_04753_),
    .A1(\u_rf.reg7_q[15] ),
    .S(_04743_),
    .X(_04754_));
 sky130_fd_sc_hd__clkbuf_1 _09917_ (.A(_04754_),
    .X(_00239_));
 sky130_fd_sc_hd__buf_2 _09918_ (.A(\u_decod.rf_ff_res_data_i[16] ),
    .X(_04755_));
 sky130_fd_sc_hd__mux2_1 _09919_ (.A0(_04755_),
    .A1(\u_rf.reg7_q[16] ),
    .S(_04743_),
    .X(_04756_));
 sky130_fd_sc_hd__clkbuf_1 _09920_ (.A(_04756_),
    .X(_00240_));
 sky130_fd_sc_hd__clkbuf_2 _09921_ (.A(\u_decod.rf_ff_res_data_i[17] ),
    .X(_04757_));
 sky130_fd_sc_hd__mux2_1 _09922_ (.A0(_04757_),
    .A1(\u_rf.reg7_q[17] ),
    .S(_04743_),
    .X(_04758_));
 sky130_fd_sc_hd__clkbuf_1 _09923_ (.A(_04758_),
    .X(_00241_));
 sky130_fd_sc_hd__clkbuf_2 _09924_ (.A(\u_decod.rf_ff_res_data_i[18] ),
    .X(_04759_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(_04759_),
    .A1(\u_rf.reg7_q[18] ),
    .S(_04743_),
    .X(_04760_));
 sky130_fd_sc_hd__clkbuf_1 _09926_ (.A(_04760_),
    .X(_00242_));
 sky130_fd_sc_hd__clkbuf_2 _09927_ (.A(\u_decod.rf_ff_res_data_i[19] ),
    .X(_04761_));
 sky130_fd_sc_hd__mux2_1 _09928_ (.A0(_04761_),
    .A1(\u_rf.reg7_q[19] ),
    .S(_04743_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_1 _09929_ (.A(_04762_),
    .X(_00243_));
 sky130_fd_sc_hd__buf_2 _09930_ (.A(\u_decod.rf_ff_res_data_i[20] ),
    .X(_04763_));
 sky130_fd_sc_hd__buf_6 _09931_ (.A(_04721_),
    .X(_04764_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(_04763_),
    .A1(\u_rf.reg7_q[20] ),
    .S(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__clkbuf_1 _09933_ (.A(_04765_),
    .X(_00244_));
 sky130_fd_sc_hd__buf_2 _09934_ (.A(\u_decod.rf_ff_res_data_i[21] ),
    .X(_04766_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(_04766_),
    .A1(\u_rf.reg7_q[21] ),
    .S(_04764_),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_1 _09936_ (.A(_04767_),
    .X(_00245_));
 sky130_fd_sc_hd__buf_2 _09937_ (.A(\u_decod.rf_ff_res_data_i[22] ),
    .X(_04768_));
 sky130_fd_sc_hd__mux2_1 _09938_ (.A0(_04768_),
    .A1(\u_rf.reg7_q[22] ),
    .S(_04764_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_1 _09939_ (.A(_04769_),
    .X(_00246_));
 sky130_fd_sc_hd__clkbuf_2 _09940_ (.A(\u_decod.rf_ff_res_data_i[23] ),
    .X(_04770_));
 sky130_fd_sc_hd__mux2_1 _09941_ (.A0(_04770_),
    .A1(\u_rf.reg7_q[23] ),
    .S(_04764_),
    .X(_04771_));
 sky130_fd_sc_hd__clkbuf_1 _09942_ (.A(_04771_),
    .X(_00247_));
 sky130_fd_sc_hd__buf_2 _09943_ (.A(\u_decod.rf_ff_res_data_i[24] ),
    .X(_04772_));
 sky130_fd_sc_hd__mux2_1 _09944_ (.A0(_04772_),
    .A1(\u_rf.reg7_q[24] ),
    .S(_04764_),
    .X(_04773_));
 sky130_fd_sc_hd__clkbuf_1 _09945_ (.A(_04773_),
    .X(_00248_));
 sky130_fd_sc_hd__buf_2 _09946_ (.A(\u_decod.rf_ff_res_data_i[25] ),
    .X(_04774_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(_04774_),
    .A1(\u_rf.reg7_q[25] ),
    .S(_04764_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_1 _09948_ (.A(_04775_),
    .X(_00249_));
 sky130_fd_sc_hd__buf_2 _09949_ (.A(\u_decod.rf_ff_res_data_i[26] ),
    .X(_04776_));
 sky130_fd_sc_hd__mux2_1 _09950_ (.A0(_04776_),
    .A1(\u_rf.reg7_q[26] ),
    .S(_04764_),
    .X(_04777_));
 sky130_fd_sc_hd__clkbuf_1 _09951_ (.A(_04777_),
    .X(_00250_));
 sky130_fd_sc_hd__clkbuf_2 _09952_ (.A(\u_decod.rf_ff_res_data_i[27] ),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(_04778_),
    .A1(\u_rf.reg7_q[27] ),
    .S(_04764_),
    .X(_04779_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_04779_),
    .X(_00251_));
 sky130_fd_sc_hd__clkbuf_2 _09955_ (.A(\u_decod.rf_ff_res_data_i[28] ),
    .X(_04780_));
 sky130_fd_sc_hd__mux2_1 _09956_ (.A0(_04780_),
    .A1(\u_rf.reg7_q[28] ),
    .S(_04764_),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_1 _09957_ (.A(_04781_),
    .X(_00252_));
 sky130_fd_sc_hd__clkbuf_2 _09958_ (.A(\u_decod.rf_ff_res_data_i[29] ),
    .X(_04782_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(_04782_),
    .A1(\u_rf.reg7_q[29] ),
    .S(_04764_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_1 _09960_ (.A(_04783_),
    .X(_00253_));
 sky130_fd_sc_hd__clkbuf_2 _09961_ (.A(\u_decod.rf_ff_res_data_i[30] ),
    .X(_04784_));
 sky130_fd_sc_hd__mux2_1 _09962_ (.A0(_04784_),
    .A1(\u_rf.reg7_q[30] ),
    .S(_04721_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_1 _09963_ (.A(_04785_),
    .X(_00254_));
 sky130_fd_sc_hd__clkbuf_2 _09964_ (.A(\u_decod.rf_ff_res_data_i[31] ),
    .X(_04786_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(_04786_),
    .A1(\u_rf.reg7_q[31] ),
    .S(_04721_),
    .X(_04787_));
 sky130_fd_sc_hd__clkbuf_1 _09966_ (.A(_04787_),
    .X(_00255_));
 sky130_fd_sc_hd__or4_4 _09967_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_04424_),
    .C(_01531_),
    .D(_01535_),
    .X(_04788_));
 sky130_fd_sc_hd__nor2_4 _09968_ (.A(_04423_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__clkbuf_8 _09969_ (.A(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__mux2_1 _09970_ (.A0(\u_rf.reg8_q[0] ),
    .A1(_04421_),
    .S(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__clkbuf_1 _09971_ (.A(_04791_),
    .X(_00256_));
 sky130_fd_sc_hd__mux2_1 _09972_ (.A0(\u_rf.reg8_q[1] ),
    .A1(_04430_),
    .S(_04790_),
    .X(_04792_));
 sky130_fd_sc_hd__clkbuf_1 _09973_ (.A(_04792_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _09974_ (.A0(\u_rf.reg8_q[2] ),
    .A1(_04432_),
    .S(_04790_),
    .X(_04793_));
 sky130_fd_sc_hd__clkbuf_1 _09975_ (.A(_04793_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _09976_ (.A0(\u_rf.reg8_q[3] ),
    .A1(_04434_),
    .S(_04790_),
    .X(_04794_));
 sky130_fd_sc_hd__clkbuf_1 _09977_ (.A(_04794_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _09978_ (.A0(\u_rf.reg8_q[4] ),
    .A1(_04436_),
    .S(_04790_),
    .X(_04795_));
 sky130_fd_sc_hd__clkbuf_1 _09979_ (.A(_04795_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _09980_ (.A0(\u_rf.reg8_q[5] ),
    .A1(_04438_),
    .S(_04790_),
    .X(_04796_));
 sky130_fd_sc_hd__clkbuf_1 _09981_ (.A(_04796_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _09982_ (.A0(\u_rf.reg8_q[6] ),
    .A1(_04440_),
    .S(_04790_),
    .X(_04797_));
 sky130_fd_sc_hd__clkbuf_1 _09983_ (.A(_04797_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _09984_ (.A0(\u_rf.reg8_q[7] ),
    .A1(_04442_),
    .S(_04790_),
    .X(_04798_));
 sky130_fd_sc_hd__clkbuf_1 _09985_ (.A(_04798_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _09986_ (.A0(\u_rf.reg8_q[8] ),
    .A1(_04444_),
    .S(_04790_),
    .X(_04799_));
 sky130_fd_sc_hd__clkbuf_1 _09987_ (.A(_04799_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _09988_ (.A0(\u_rf.reg8_q[9] ),
    .A1(_04446_),
    .S(_04790_),
    .X(_04800_));
 sky130_fd_sc_hd__clkbuf_1 _09989_ (.A(_04800_),
    .X(_00265_));
 sky130_fd_sc_hd__buf_6 _09990_ (.A(_04789_),
    .X(_04801_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(\u_rf.reg8_q[10] ),
    .A1(_04448_),
    .S(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__clkbuf_1 _09992_ (.A(_04802_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _09993_ (.A0(\u_rf.reg8_q[11] ),
    .A1(_04451_),
    .S(_04801_),
    .X(_04803_));
 sky130_fd_sc_hd__clkbuf_1 _09994_ (.A(_04803_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(\u_rf.reg8_q[12] ),
    .A1(_04453_),
    .S(_04801_),
    .X(_04804_));
 sky130_fd_sc_hd__clkbuf_1 _09996_ (.A(_04804_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _09997_ (.A0(\u_rf.reg8_q[13] ),
    .A1(_04455_),
    .S(_04801_),
    .X(_04805_));
 sky130_fd_sc_hd__clkbuf_1 _09998_ (.A(_04805_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(\u_rf.reg8_q[14] ),
    .A1(_04457_),
    .S(_04801_),
    .X(_04806_));
 sky130_fd_sc_hd__clkbuf_1 _10000_ (.A(_04806_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(\u_rf.reg8_q[15] ),
    .A1(_04459_),
    .S(_04801_),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_1 _10002_ (.A(_04807_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(\u_rf.reg8_q[16] ),
    .A1(_04461_),
    .S(_04801_),
    .X(_04808_));
 sky130_fd_sc_hd__clkbuf_1 _10004_ (.A(_04808_),
    .X(_00272_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(\u_rf.reg8_q[17] ),
    .A1(_04463_),
    .S(_04801_),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_1 _10006_ (.A(_04809_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(\u_rf.reg8_q[18] ),
    .A1(_04465_),
    .S(_04801_),
    .X(_04810_));
 sky130_fd_sc_hd__clkbuf_1 _10008_ (.A(_04810_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(\u_rf.reg8_q[19] ),
    .A1(_04467_),
    .S(_04801_),
    .X(_04811_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_04811_),
    .X(_00275_));
 sky130_fd_sc_hd__clkbuf_8 _10011_ (.A(_04789_),
    .X(_04812_));
 sky130_fd_sc_hd__mux2_1 _10012_ (.A0(\u_rf.reg8_q[20] ),
    .A1(_04469_),
    .S(_04812_),
    .X(_04813_));
 sky130_fd_sc_hd__clkbuf_1 _10013_ (.A(_04813_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _10014_ (.A0(\u_rf.reg8_q[21] ),
    .A1(_04472_),
    .S(_04812_),
    .X(_04814_));
 sky130_fd_sc_hd__clkbuf_1 _10015_ (.A(_04814_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _10016_ (.A0(\u_rf.reg8_q[22] ),
    .A1(_04474_),
    .S(_04812_),
    .X(_04815_));
 sky130_fd_sc_hd__clkbuf_1 _10017_ (.A(_04815_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _10018_ (.A0(\u_rf.reg8_q[23] ),
    .A1(_04476_),
    .S(_04812_),
    .X(_04816_));
 sky130_fd_sc_hd__clkbuf_1 _10019_ (.A(_04816_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _10020_ (.A0(\u_rf.reg8_q[24] ),
    .A1(_04478_),
    .S(_04812_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _10021_ (.A(_04817_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _10022_ (.A0(\u_rf.reg8_q[25] ),
    .A1(_04480_),
    .S(_04812_),
    .X(_04818_));
 sky130_fd_sc_hd__clkbuf_1 _10023_ (.A(_04818_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _10024_ (.A0(\u_rf.reg8_q[26] ),
    .A1(_04482_),
    .S(_04812_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _10025_ (.A(_04819_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _10026_ (.A0(\u_rf.reg8_q[27] ),
    .A1(_04484_),
    .S(_04812_),
    .X(_04820_));
 sky130_fd_sc_hd__clkbuf_1 _10027_ (.A(_04820_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _10028_ (.A0(\u_rf.reg8_q[28] ),
    .A1(_04486_),
    .S(_04812_),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_1 _10029_ (.A(_04821_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _10030_ (.A0(\u_rf.reg8_q[29] ),
    .A1(_04488_),
    .S(_04812_),
    .X(_04822_));
 sky130_fd_sc_hd__clkbuf_1 _10031_ (.A(_04822_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _10032_ (.A0(\u_rf.reg8_q[30] ),
    .A1(_04490_),
    .S(_04789_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_1 _10033_ (.A(_04823_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _10034_ (.A0(\u_rf.reg8_q[31] ),
    .A1(_04492_),
    .S(_04789_),
    .X(_04824_));
 sky130_fd_sc_hd__clkbuf_1 _10035_ (.A(_04824_),
    .X(_00287_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(_01531_),
    .B(_01535_),
    .Y(_04825_));
 sky130_fd_sc_hd__and3_4 _10037_ (.A(_04643_),
    .B(_04644_),
    .C(_04825_),
    .X(_04826_));
 sky130_fd_sc_hd__buf_4 _10038_ (.A(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(\u_rf.reg9_q[0] ),
    .A1(_04421_),
    .S(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__clkbuf_1 _10040_ (.A(_04828_),
    .X(_00288_));
 sky130_fd_sc_hd__mux2_1 _10041_ (.A0(\u_rf.reg9_q[1] ),
    .A1(_04430_),
    .S(_04827_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _10042_ (.A(_04829_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(\u_rf.reg9_q[2] ),
    .A1(_04432_),
    .S(_04827_),
    .X(_04830_));
 sky130_fd_sc_hd__clkbuf_1 _10044_ (.A(_04830_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(\u_rf.reg9_q[3] ),
    .A1(_04434_),
    .S(_04827_),
    .X(_04831_));
 sky130_fd_sc_hd__clkbuf_1 _10046_ (.A(_04831_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(\u_rf.reg9_q[4] ),
    .A1(_04436_),
    .S(_04827_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_1 _10048_ (.A(_04832_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(\u_rf.reg9_q[5] ),
    .A1(_04438_),
    .S(_04827_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _10050_ (.A(_04833_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _10051_ (.A0(\u_rf.reg9_q[6] ),
    .A1(_04440_),
    .S(_04827_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_1 _10052_ (.A(_04834_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(\u_rf.reg9_q[7] ),
    .A1(_04442_),
    .S(_04827_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _10054_ (.A(_04835_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(\u_rf.reg9_q[8] ),
    .A1(_04444_),
    .S(_04827_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _10056_ (.A(_04836_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _10057_ (.A0(\u_rf.reg9_q[9] ),
    .A1(_04446_),
    .S(_04827_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _10058_ (.A(_04837_),
    .X(_00297_));
 sky130_fd_sc_hd__buf_8 _10059_ (.A(_04826_),
    .X(_04838_));
 sky130_fd_sc_hd__mux2_1 _10060_ (.A0(\u_rf.reg9_q[10] ),
    .A1(_04448_),
    .S(_04838_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _10061_ (.A(_04839_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(\u_rf.reg9_q[11] ),
    .A1(_04451_),
    .S(_04838_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _10063_ (.A(_04840_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(\u_rf.reg9_q[12] ),
    .A1(_04453_),
    .S(_04838_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _10065_ (.A(_04841_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(\u_rf.reg9_q[13] ),
    .A1(_04455_),
    .S(_04838_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _10067_ (.A(_04842_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(\u_rf.reg9_q[14] ),
    .A1(_04457_),
    .S(_04838_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _10069_ (.A(_04843_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _10070_ (.A0(\u_rf.reg9_q[15] ),
    .A1(_04459_),
    .S(_04838_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _10071_ (.A(_04844_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _10072_ (.A0(\u_rf.reg9_q[16] ),
    .A1(_04461_),
    .S(_04838_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _10073_ (.A(_04845_),
    .X(_00304_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(\u_rf.reg9_q[17] ),
    .A1(_04463_),
    .S(_04838_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _10075_ (.A(_04846_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(\u_rf.reg9_q[18] ),
    .A1(_04465_),
    .S(_04838_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _10077_ (.A(_04847_),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(\u_rf.reg9_q[19] ),
    .A1(_04467_),
    .S(_04838_),
    .X(_04848_));
 sky130_fd_sc_hd__clkbuf_1 _10079_ (.A(_04848_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_4 _10080_ (.A(_04826_),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_1 _10081_ (.A0(\u_rf.reg9_q[20] ),
    .A1(_04469_),
    .S(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__clkbuf_1 _10082_ (.A(_04850_),
    .X(_00308_));
 sky130_fd_sc_hd__mux2_1 _10083_ (.A0(\u_rf.reg9_q[21] ),
    .A1(_04472_),
    .S(_04849_),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_1 _10084_ (.A(_04851_),
    .X(_00309_));
 sky130_fd_sc_hd__mux2_1 _10085_ (.A0(\u_rf.reg9_q[22] ),
    .A1(_04474_),
    .S(_04849_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _10086_ (.A(_04852_),
    .X(_00310_));
 sky130_fd_sc_hd__mux2_1 _10087_ (.A0(\u_rf.reg9_q[23] ),
    .A1(_04476_),
    .S(_04849_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _10088_ (.A(_04853_),
    .X(_00311_));
 sky130_fd_sc_hd__mux2_1 _10089_ (.A0(\u_rf.reg9_q[24] ),
    .A1(_04478_),
    .S(_04849_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _10090_ (.A(_04854_),
    .X(_00312_));
 sky130_fd_sc_hd__mux2_1 _10091_ (.A0(\u_rf.reg9_q[25] ),
    .A1(_04480_),
    .S(_04849_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _10092_ (.A(_04855_),
    .X(_00313_));
 sky130_fd_sc_hd__mux2_1 _10093_ (.A0(\u_rf.reg9_q[26] ),
    .A1(_04482_),
    .S(_04849_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_1 _10094_ (.A(_04856_),
    .X(_00314_));
 sky130_fd_sc_hd__mux2_1 _10095_ (.A0(\u_rf.reg9_q[27] ),
    .A1(_04484_),
    .S(_04849_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _10096_ (.A(_04857_),
    .X(_00315_));
 sky130_fd_sc_hd__mux2_1 _10097_ (.A0(\u_rf.reg9_q[28] ),
    .A1(_04486_),
    .S(_04849_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _10098_ (.A(_04858_),
    .X(_00316_));
 sky130_fd_sc_hd__mux2_1 _10099_ (.A0(\u_rf.reg9_q[29] ),
    .A1(_04488_),
    .S(_04849_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _10100_ (.A(_04859_),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _10101_ (.A0(\u_rf.reg9_q[30] ),
    .A1(_04490_),
    .S(_04826_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _10102_ (.A(_04860_),
    .X(_00318_));
 sky130_fd_sc_hd__mux2_1 _10103_ (.A0(\u_rf.reg9_q[31] ),
    .A1(_04492_),
    .S(_04826_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _10104_ (.A(_04861_),
    .X(_00319_));
 sky130_fd_sc_hd__and3_2 _10105_ (.A(_04643_),
    .B(_04682_),
    .C(_04825_),
    .X(_04862_));
 sky130_fd_sc_hd__buf_6 _10106_ (.A(_04862_),
    .X(_04863_));
 sky130_fd_sc_hd__mux2_1 _10107_ (.A0(\u_rf.reg10_q[0] ),
    .A1(_04421_),
    .S(_04863_),
    .X(_04864_));
 sky130_fd_sc_hd__clkbuf_1 _10108_ (.A(_04864_),
    .X(_00320_));
 sky130_fd_sc_hd__mux2_1 _10109_ (.A0(\u_rf.reg10_q[1] ),
    .A1(_04430_),
    .S(_04863_),
    .X(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _10110_ (.A(_04865_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _10111_ (.A0(\u_rf.reg10_q[2] ),
    .A1(_04432_),
    .S(_04863_),
    .X(_04866_));
 sky130_fd_sc_hd__clkbuf_1 _10112_ (.A(_04866_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _10113_ (.A0(\u_rf.reg10_q[3] ),
    .A1(_04434_),
    .S(_04863_),
    .X(_04867_));
 sky130_fd_sc_hd__clkbuf_1 _10114_ (.A(_04867_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _10115_ (.A0(\u_rf.reg10_q[4] ),
    .A1(_04436_),
    .S(_04863_),
    .X(_04868_));
 sky130_fd_sc_hd__clkbuf_1 _10116_ (.A(_04868_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _10117_ (.A0(\u_rf.reg10_q[5] ),
    .A1(_04438_),
    .S(_04863_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _10118_ (.A(_04869_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _10119_ (.A0(\u_rf.reg10_q[6] ),
    .A1(_04440_),
    .S(_04863_),
    .X(_04870_));
 sky130_fd_sc_hd__clkbuf_1 _10120_ (.A(_04870_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _10121_ (.A0(\u_rf.reg10_q[7] ),
    .A1(_04442_),
    .S(_04863_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _10122_ (.A(_04871_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _10123_ (.A0(\u_rf.reg10_q[8] ),
    .A1(_04444_),
    .S(_04863_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _10124_ (.A(_04872_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _10125_ (.A0(\u_rf.reg10_q[9] ),
    .A1(_04446_),
    .S(_04863_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _10126_ (.A(_04873_),
    .X(_00329_));
 sky130_fd_sc_hd__buf_6 _10127_ (.A(_04862_),
    .X(_04874_));
 sky130_fd_sc_hd__mux2_1 _10128_ (.A0(\u_rf.reg10_q[10] ),
    .A1(_04448_),
    .S(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_1 _10129_ (.A(_04875_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(\u_rf.reg10_q[11] ),
    .A1(_04451_),
    .S(_04874_),
    .X(_04876_));
 sky130_fd_sc_hd__clkbuf_1 _10131_ (.A(_04876_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _10132_ (.A0(\u_rf.reg10_q[12] ),
    .A1(_04453_),
    .S(_04874_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _10133_ (.A(_04877_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _10134_ (.A0(\u_rf.reg10_q[13] ),
    .A1(_04455_),
    .S(_04874_),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_1 _10135_ (.A(_04878_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(\u_rf.reg10_q[14] ),
    .A1(_04457_),
    .S(_04874_),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _10137_ (.A(_04879_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _10138_ (.A0(\u_rf.reg10_q[15] ),
    .A1(_04459_),
    .S(_04874_),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _10139_ (.A(_04880_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _10140_ (.A0(\u_rf.reg10_q[16] ),
    .A1(_04461_),
    .S(_04874_),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _10141_ (.A(_04881_),
    .X(_00336_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(\u_rf.reg10_q[17] ),
    .A1(_04463_),
    .S(_04874_),
    .X(_04882_));
 sky130_fd_sc_hd__clkbuf_1 _10143_ (.A(_04882_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _10144_ (.A0(\u_rf.reg10_q[18] ),
    .A1(_04465_),
    .S(_04874_),
    .X(_04883_));
 sky130_fd_sc_hd__clkbuf_1 _10145_ (.A(_04883_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _10146_ (.A0(\u_rf.reg10_q[19] ),
    .A1(_04467_),
    .S(_04874_),
    .X(_04884_));
 sky130_fd_sc_hd__clkbuf_1 _10147_ (.A(_04884_),
    .X(_00339_));
 sky130_fd_sc_hd__clkbuf_8 _10148_ (.A(_04862_),
    .X(_04885_));
 sky130_fd_sc_hd__mux2_1 _10149_ (.A0(\u_rf.reg10_q[20] ),
    .A1(_04469_),
    .S(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__clkbuf_1 _10150_ (.A(_04886_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(\u_rf.reg10_q[21] ),
    .A1(_04472_),
    .S(_04885_),
    .X(_04887_));
 sky130_fd_sc_hd__clkbuf_1 _10152_ (.A(_04887_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _10153_ (.A0(\u_rf.reg10_q[22] ),
    .A1(_04474_),
    .S(_04885_),
    .X(_04888_));
 sky130_fd_sc_hd__clkbuf_1 _10154_ (.A(_04888_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _10155_ (.A0(\u_rf.reg10_q[23] ),
    .A1(_04476_),
    .S(_04885_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_1 _10156_ (.A(_04889_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(\u_rf.reg10_q[24] ),
    .A1(_04478_),
    .S(_04885_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_1 _10158_ (.A(_04890_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _10159_ (.A0(\u_rf.reg10_q[25] ),
    .A1(_04480_),
    .S(_04885_),
    .X(_04891_));
 sky130_fd_sc_hd__clkbuf_1 _10160_ (.A(_04891_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(\u_rf.reg10_q[26] ),
    .A1(_04482_),
    .S(_04885_),
    .X(_04892_));
 sky130_fd_sc_hd__clkbuf_1 _10162_ (.A(_04892_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(\u_rf.reg10_q[27] ),
    .A1(_04484_),
    .S(_04885_),
    .X(_04893_));
 sky130_fd_sc_hd__clkbuf_1 _10164_ (.A(_04893_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _10165_ (.A0(\u_rf.reg10_q[28] ),
    .A1(_04486_),
    .S(_04885_),
    .X(_04894_));
 sky130_fd_sc_hd__clkbuf_1 _10166_ (.A(_04894_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _10167_ (.A0(\u_rf.reg10_q[29] ),
    .A1(_04488_),
    .S(_04885_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_1 _10168_ (.A(_04895_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(\u_rf.reg10_q[30] ),
    .A1(_04490_),
    .S(_04862_),
    .X(_04896_));
 sky130_fd_sc_hd__clkbuf_1 _10170_ (.A(_04896_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(\u_rf.reg10_q[31] ),
    .A1(_04492_),
    .S(_04862_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_1 _10172_ (.A(_04897_),
    .X(_00351_));
 sky130_fd_sc_hd__or3b_1 _10173_ (.A(_04422_),
    .B(_04568_),
    .C_N(_04825_),
    .X(_04898_));
 sky130_fd_sc_hd__buf_2 _10174_ (.A(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_8 _10175_ (.A(_04899_),
    .X(_04900_));
 sky130_fd_sc_hd__mux2_1 _10176_ (.A0(_04719_),
    .A1(\u_rf.reg11_q[0] ),
    .S(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_1 _10177_ (.A(_04901_),
    .X(_00352_));
 sky130_fd_sc_hd__mux2_1 _10178_ (.A0(_04724_),
    .A1(\u_rf.reg11_q[1] ),
    .S(_04900_),
    .X(_04902_));
 sky130_fd_sc_hd__clkbuf_1 _10179_ (.A(_04902_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(_04726_),
    .A1(\u_rf.reg11_q[2] ),
    .S(_04900_),
    .X(_04903_));
 sky130_fd_sc_hd__clkbuf_1 _10181_ (.A(_04903_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(_04728_),
    .A1(\u_rf.reg11_q[3] ),
    .S(_04900_),
    .X(_04904_));
 sky130_fd_sc_hd__clkbuf_1 _10183_ (.A(_04904_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(_04730_),
    .A1(\u_rf.reg11_q[4] ),
    .S(_04900_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_1 _10185_ (.A(_04905_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(_04732_),
    .A1(\u_rf.reg11_q[5] ),
    .S(_04900_),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_1 _10187_ (.A(_04906_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(_04734_),
    .A1(\u_rf.reg11_q[6] ),
    .S(_04900_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_1 _10189_ (.A(_04907_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(_04736_),
    .A1(\u_rf.reg11_q[7] ),
    .S(_04900_),
    .X(_04908_));
 sky130_fd_sc_hd__clkbuf_1 _10191_ (.A(_04908_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(_04738_),
    .A1(\u_rf.reg11_q[8] ),
    .S(_04900_),
    .X(_04909_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_04909_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(_04740_),
    .A1(\u_rf.reg11_q[9] ),
    .S(_04900_),
    .X(_04910_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_04910_),
    .X(_00361_));
 sky130_fd_sc_hd__buf_6 _10196_ (.A(_04899_),
    .X(_04911_));
 sky130_fd_sc_hd__mux2_1 _10197_ (.A0(_04742_),
    .A1(\u_rf.reg11_q[10] ),
    .S(_04911_),
    .X(_04912_));
 sky130_fd_sc_hd__clkbuf_1 _10198_ (.A(_04912_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(_04745_),
    .A1(\u_rf.reg11_q[11] ),
    .S(_04911_),
    .X(_04913_));
 sky130_fd_sc_hd__clkbuf_1 _10200_ (.A(_04913_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(_04747_),
    .A1(\u_rf.reg11_q[12] ),
    .S(_04911_),
    .X(_04914_));
 sky130_fd_sc_hd__clkbuf_1 _10202_ (.A(_04914_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(_04749_),
    .A1(\u_rf.reg11_q[13] ),
    .S(_04911_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_1 _10204_ (.A(_04915_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _10205_ (.A0(_04751_),
    .A1(\u_rf.reg11_q[14] ),
    .S(_04911_),
    .X(_04916_));
 sky130_fd_sc_hd__clkbuf_1 _10206_ (.A(_04916_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _10207_ (.A0(_04753_),
    .A1(\u_rf.reg11_q[15] ),
    .S(_04911_),
    .X(_04917_));
 sky130_fd_sc_hd__clkbuf_1 _10208_ (.A(_04917_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _10209_ (.A0(_04755_),
    .A1(\u_rf.reg11_q[16] ),
    .S(_04911_),
    .X(_04918_));
 sky130_fd_sc_hd__clkbuf_1 _10210_ (.A(_04918_),
    .X(_00368_));
 sky130_fd_sc_hd__mux2_1 _10211_ (.A0(_04757_),
    .A1(\u_rf.reg11_q[17] ),
    .S(_04911_),
    .X(_04919_));
 sky130_fd_sc_hd__clkbuf_1 _10212_ (.A(_04919_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _10213_ (.A0(_04759_),
    .A1(\u_rf.reg11_q[18] ),
    .S(_04911_),
    .X(_04920_));
 sky130_fd_sc_hd__clkbuf_1 _10214_ (.A(_04920_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(_04761_),
    .A1(\u_rf.reg11_q[19] ),
    .S(_04911_),
    .X(_04921_));
 sky130_fd_sc_hd__clkbuf_1 _10216_ (.A(_04921_),
    .X(_00371_));
 sky130_fd_sc_hd__clkbuf_8 _10217_ (.A(_04899_),
    .X(_04922_));
 sky130_fd_sc_hd__mux2_1 _10218_ (.A0(_04763_),
    .A1(\u_rf.reg11_q[20] ),
    .S(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_1 _10219_ (.A(_04923_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _10220_ (.A0(_04766_),
    .A1(\u_rf.reg11_q[21] ),
    .S(_04922_),
    .X(_04924_));
 sky130_fd_sc_hd__clkbuf_1 _10221_ (.A(_04924_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _10222_ (.A0(_04768_),
    .A1(\u_rf.reg11_q[22] ),
    .S(_04922_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_1 _10223_ (.A(_04925_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _10224_ (.A0(_04770_),
    .A1(\u_rf.reg11_q[23] ),
    .S(_04922_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _10225_ (.A(_04926_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _10226_ (.A0(_04772_),
    .A1(\u_rf.reg11_q[24] ),
    .S(_04922_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_1 _10227_ (.A(_04927_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _10228_ (.A0(_04774_),
    .A1(\u_rf.reg11_q[25] ),
    .S(_04922_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _10229_ (.A(_04928_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _10230_ (.A0(_04776_),
    .A1(\u_rf.reg11_q[26] ),
    .S(_04922_),
    .X(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _10231_ (.A(_04929_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _10232_ (.A0(_04778_),
    .A1(\u_rf.reg11_q[27] ),
    .S(_04922_),
    .X(_04930_));
 sky130_fd_sc_hd__clkbuf_1 _10233_ (.A(_04930_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _10234_ (.A0(_04780_),
    .A1(\u_rf.reg11_q[28] ),
    .S(_04922_),
    .X(_04931_));
 sky130_fd_sc_hd__clkbuf_1 _10235_ (.A(_04931_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _10236_ (.A0(_04782_),
    .A1(\u_rf.reg11_q[29] ),
    .S(_04922_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _10237_ (.A(_04932_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _10238_ (.A0(_04784_),
    .A1(\u_rf.reg11_q[30] ),
    .S(_04899_),
    .X(_04933_));
 sky130_fd_sc_hd__clkbuf_1 _10239_ (.A(_04933_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _10240_ (.A0(_04786_),
    .A1(\u_rf.reg11_q[31] ),
    .S(_04899_),
    .X(_04934_));
 sky130_fd_sc_hd__clkbuf_1 _10241_ (.A(_04934_),
    .X(_00383_));
 sky130_fd_sc_hd__buf_2 _10242_ (.A(\u_decod.rf_ff_res_data_i[0] ),
    .X(_04935_));
 sky130_fd_sc_hd__nand2_2 _10243_ (.A(_01531_),
    .B(_01536_),
    .Y(_04936_));
 sky130_fd_sc_hd__or3_2 _10244_ (.A(\u_decod.rf_ff_rd_adr_q_i[0] ),
    .B(_04424_),
    .C(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_2 _10245_ (.A(_04423_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__clkbuf_8 _10246_ (.A(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__mux2_1 _10247_ (.A0(\u_rf.reg12_q[0] ),
    .A1(_04935_),
    .S(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_1 _10248_ (.A(_04940_),
    .X(_00384_));
 sky130_fd_sc_hd__clkbuf_2 _10249_ (.A(\u_decod.rf_ff_res_data_i[1] ),
    .X(_04941_));
 sky130_fd_sc_hd__mux2_1 _10250_ (.A0(\u_rf.reg12_q[1] ),
    .A1(_04941_),
    .S(_04939_),
    .X(_04942_));
 sky130_fd_sc_hd__clkbuf_1 _10251_ (.A(_04942_),
    .X(_00385_));
 sky130_fd_sc_hd__buf_2 _10252_ (.A(\u_decod.rf_ff_res_data_i[2] ),
    .X(_04943_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(\u_rf.reg12_q[2] ),
    .A1(_04943_),
    .S(_04939_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_1 _10254_ (.A(_04944_),
    .X(_00386_));
 sky130_fd_sc_hd__buf_2 _10255_ (.A(\u_decod.rf_ff_res_data_i[3] ),
    .X(_04945_));
 sky130_fd_sc_hd__mux2_1 _10256_ (.A0(\u_rf.reg12_q[3] ),
    .A1(_04945_),
    .S(_04939_),
    .X(_04946_));
 sky130_fd_sc_hd__clkbuf_1 _10257_ (.A(_04946_),
    .X(_00387_));
 sky130_fd_sc_hd__clkbuf_2 _10258_ (.A(\u_decod.rf_ff_res_data_i[4] ),
    .X(_04947_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(\u_rf.reg12_q[4] ),
    .A1(_04947_),
    .S(_04939_),
    .X(_04948_));
 sky130_fd_sc_hd__clkbuf_1 _10260_ (.A(_04948_),
    .X(_00388_));
 sky130_fd_sc_hd__buf_2 _10261_ (.A(\u_decod.rf_ff_res_data_i[5] ),
    .X(_04949_));
 sky130_fd_sc_hd__mux2_1 _10262_ (.A0(\u_rf.reg12_q[5] ),
    .A1(_04949_),
    .S(_04939_),
    .X(_04950_));
 sky130_fd_sc_hd__clkbuf_1 _10263_ (.A(_04950_),
    .X(_00389_));
 sky130_fd_sc_hd__buf_2 _10264_ (.A(\u_decod.rf_ff_res_data_i[6] ),
    .X(_04951_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(\u_rf.reg12_q[6] ),
    .A1(_04951_),
    .S(_04939_),
    .X(_04952_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_04952_),
    .X(_00390_));
 sky130_fd_sc_hd__clkbuf_2 _10267_ (.A(\u_decod.rf_ff_res_data_i[7] ),
    .X(_04953_));
 sky130_fd_sc_hd__mux2_1 _10268_ (.A0(\u_rf.reg12_q[7] ),
    .A1(_04953_),
    .S(_04939_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_1 _10269_ (.A(_04954_),
    .X(_00391_));
 sky130_fd_sc_hd__clkbuf_2 _10270_ (.A(\u_decod.rf_ff_res_data_i[8] ),
    .X(_04955_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(\u_rf.reg12_q[8] ),
    .A1(_04955_),
    .S(_04939_),
    .X(_04956_));
 sky130_fd_sc_hd__clkbuf_1 _10272_ (.A(_04956_),
    .X(_00392_));
 sky130_fd_sc_hd__buf_2 _10273_ (.A(\u_decod.rf_ff_res_data_i[9] ),
    .X(_04957_));
 sky130_fd_sc_hd__mux2_1 _10274_ (.A0(\u_rf.reg12_q[9] ),
    .A1(_04957_),
    .S(_04939_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_1 _10275_ (.A(_04958_),
    .X(_00393_));
 sky130_fd_sc_hd__buf_2 _10276_ (.A(\u_decod.rf_ff_res_data_i[10] ),
    .X(_04959_));
 sky130_fd_sc_hd__clkbuf_8 _10277_ (.A(_04938_),
    .X(_04960_));
 sky130_fd_sc_hd__mux2_1 _10278_ (.A0(\u_rf.reg12_q[10] ),
    .A1(_04959_),
    .S(_04960_),
    .X(_04961_));
 sky130_fd_sc_hd__clkbuf_1 _10279_ (.A(_04961_),
    .X(_00394_));
 sky130_fd_sc_hd__clkbuf_2 _10280_ (.A(\u_decod.rf_ff_res_data_i[11] ),
    .X(_04962_));
 sky130_fd_sc_hd__mux2_1 _10281_ (.A0(\u_rf.reg12_q[11] ),
    .A1(_04962_),
    .S(_04960_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_1 _10282_ (.A(_04963_),
    .X(_00395_));
 sky130_fd_sc_hd__clkbuf_2 _10283_ (.A(\u_decod.rf_ff_res_data_i[12] ),
    .X(_04964_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(\u_rf.reg12_q[12] ),
    .A1(_04964_),
    .S(_04960_),
    .X(_04965_));
 sky130_fd_sc_hd__clkbuf_1 _10285_ (.A(_04965_),
    .X(_00396_));
 sky130_fd_sc_hd__buf_2 _10286_ (.A(\u_decod.rf_ff_res_data_i[13] ),
    .X(_04966_));
 sky130_fd_sc_hd__mux2_1 _10287_ (.A0(\u_rf.reg12_q[13] ),
    .A1(_04966_),
    .S(_04960_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_1 _10288_ (.A(_04967_),
    .X(_00397_));
 sky130_fd_sc_hd__buf_2 _10289_ (.A(\u_decod.rf_ff_res_data_i[14] ),
    .X(_04968_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(\u_rf.reg12_q[14] ),
    .A1(_04968_),
    .S(_04960_),
    .X(_04969_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_04969_),
    .X(_00398_));
 sky130_fd_sc_hd__clkbuf_2 _10292_ (.A(\u_decod.rf_ff_res_data_i[15] ),
    .X(_04970_));
 sky130_fd_sc_hd__mux2_1 _10293_ (.A0(\u_rf.reg12_q[15] ),
    .A1(_04970_),
    .S(_04960_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_1 _10294_ (.A(_04971_),
    .X(_00399_));
 sky130_fd_sc_hd__buf_2 _10295_ (.A(\u_decod.rf_ff_res_data_i[16] ),
    .X(_04972_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(\u_rf.reg12_q[16] ),
    .A1(_04972_),
    .S(_04960_),
    .X(_04973_));
 sky130_fd_sc_hd__clkbuf_1 _10297_ (.A(_04973_),
    .X(_00400_));
 sky130_fd_sc_hd__buf_2 _10298_ (.A(\u_decod.rf_ff_res_data_i[17] ),
    .X(_04974_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(\u_rf.reg12_q[17] ),
    .A1(_04974_),
    .S(_04960_),
    .X(_04975_));
 sky130_fd_sc_hd__clkbuf_1 _10300_ (.A(_04975_),
    .X(_00401_));
 sky130_fd_sc_hd__clkbuf_2 _10301_ (.A(\u_decod.rf_ff_res_data_i[18] ),
    .X(_04976_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(\u_rf.reg12_q[18] ),
    .A1(_04976_),
    .S(_04960_),
    .X(_04977_));
 sky130_fd_sc_hd__clkbuf_1 _10303_ (.A(_04977_),
    .X(_00402_));
 sky130_fd_sc_hd__clkbuf_2 _10304_ (.A(\u_decod.rf_ff_res_data_i[19] ),
    .X(_04978_));
 sky130_fd_sc_hd__mux2_1 _10305_ (.A0(\u_rf.reg12_q[19] ),
    .A1(_04978_),
    .S(_04960_),
    .X(_04979_));
 sky130_fd_sc_hd__clkbuf_1 _10306_ (.A(_04979_),
    .X(_00403_));
 sky130_fd_sc_hd__buf_2 _10307_ (.A(\u_decod.rf_ff_res_data_i[20] ),
    .X(_04980_));
 sky130_fd_sc_hd__clkbuf_8 _10308_ (.A(_04938_),
    .X(_04981_));
 sky130_fd_sc_hd__mux2_1 _10309_ (.A0(\u_rf.reg12_q[20] ),
    .A1(_04980_),
    .S(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_1 _10310_ (.A(_04982_),
    .X(_00404_));
 sky130_fd_sc_hd__buf_2 _10311_ (.A(\u_decod.rf_ff_res_data_i[21] ),
    .X(_04983_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(\u_rf.reg12_q[21] ),
    .A1(_04983_),
    .S(_04981_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_1 _10313_ (.A(_04984_),
    .X(_00405_));
 sky130_fd_sc_hd__buf_2 _10314_ (.A(\u_decod.rf_ff_res_data_i[22] ),
    .X(_04985_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(\u_rf.reg12_q[22] ),
    .A1(_04985_),
    .S(_04981_),
    .X(_04986_));
 sky130_fd_sc_hd__clkbuf_1 _10316_ (.A(_04986_),
    .X(_00406_));
 sky130_fd_sc_hd__buf_2 _10317_ (.A(\u_decod.rf_ff_res_data_i[23] ),
    .X(_04987_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(\u_rf.reg12_q[23] ),
    .A1(_04987_),
    .S(_04981_),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_1 _10319_ (.A(_04988_),
    .X(_00407_));
 sky130_fd_sc_hd__buf_2 _10320_ (.A(\u_decod.rf_ff_res_data_i[24] ),
    .X(_04989_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(\u_rf.reg12_q[24] ),
    .A1(_04989_),
    .S(_04981_),
    .X(_04990_));
 sky130_fd_sc_hd__clkbuf_1 _10322_ (.A(_04990_),
    .X(_00408_));
 sky130_fd_sc_hd__buf_2 _10323_ (.A(\u_decod.rf_ff_res_data_i[25] ),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_1 _10324_ (.A0(\u_rf.reg12_q[25] ),
    .A1(_04991_),
    .S(_04981_),
    .X(_04992_));
 sky130_fd_sc_hd__clkbuf_1 _10325_ (.A(_04992_),
    .X(_00409_));
 sky130_fd_sc_hd__buf_2 _10326_ (.A(\u_decod.rf_ff_res_data_i[26] ),
    .X(_04993_));
 sky130_fd_sc_hd__mux2_1 _10327_ (.A0(\u_rf.reg12_q[26] ),
    .A1(_04993_),
    .S(_04981_),
    .X(_04994_));
 sky130_fd_sc_hd__clkbuf_1 _10328_ (.A(_04994_),
    .X(_00410_));
 sky130_fd_sc_hd__buf_2 _10329_ (.A(\u_decod.rf_ff_res_data_i[27] ),
    .X(_04995_));
 sky130_fd_sc_hd__mux2_1 _10330_ (.A0(\u_rf.reg12_q[27] ),
    .A1(_04995_),
    .S(_04981_),
    .X(_04996_));
 sky130_fd_sc_hd__clkbuf_1 _10331_ (.A(_04996_),
    .X(_00411_));
 sky130_fd_sc_hd__clkbuf_2 _10332_ (.A(\u_decod.rf_ff_res_data_i[28] ),
    .X(_04997_));
 sky130_fd_sc_hd__mux2_1 _10333_ (.A0(\u_rf.reg12_q[28] ),
    .A1(_04997_),
    .S(_04981_),
    .X(_04998_));
 sky130_fd_sc_hd__clkbuf_1 _10334_ (.A(_04998_),
    .X(_00412_));
 sky130_fd_sc_hd__buf_2 _10335_ (.A(\u_decod.rf_ff_res_data_i[29] ),
    .X(_04999_));
 sky130_fd_sc_hd__mux2_1 _10336_ (.A0(\u_rf.reg12_q[29] ),
    .A1(_04999_),
    .S(_04981_),
    .X(_05000_));
 sky130_fd_sc_hd__clkbuf_1 _10337_ (.A(_05000_),
    .X(_00413_));
 sky130_fd_sc_hd__buf_2 _10338_ (.A(\u_decod.rf_ff_res_data_i[30] ),
    .X(_05001_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(\u_rf.reg12_q[30] ),
    .A1(_05001_),
    .S(_04938_),
    .X(_05002_));
 sky130_fd_sc_hd__clkbuf_1 _10340_ (.A(_05002_),
    .X(_00414_));
 sky130_fd_sc_hd__buf_2 _10341_ (.A(\u_decod.rf_ff_res_data_i[31] ),
    .X(_05003_));
 sky130_fd_sc_hd__mux2_1 _10342_ (.A0(\u_rf.reg12_q[31] ),
    .A1(_05003_),
    .S(_04938_),
    .X(_05004_));
 sky130_fd_sc_hd__clkbuf_1 _10343_ (.A(_05004_),
    .X(_00415_));
 sky130_fd_sc_hd__or4_4 _10344_ (.A(_01534_),
    .B(_04424_),
    .C(_04423_),
    .D(_04936_),
    .X(_05005_));
 sky130_fd_sc_hd__buf_6 _10345_ (.A(_05005_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _10346_ (.A0(_04719_),
    .A1(\u_rf.reg13_q[0] ),
    .S(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _10347_ (.A(_05007_),
    .X(_00416_));
 sky130_fd_sc_hd__mux2_1 _10348_ (.A0(_04724_),
    .A1(\u_rf.reg13_q[1] ),
    .S(_05006_),
    .X(_05008_));
 sky130_fd_sc_hd__clkbuf_1 _10349_ (.A(_05008_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _10350_ (.A0(_04726_),
    .A1(\u_rf.reg13_q[2] ),
    .S(_05006_),
    .X(_05009_));
 sky130_fd_sc_hd__clkbuf_1 _10351_ (.A(_05009_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _10352_ (.A0(_04728_),
    .A1(\u_rf.reg13_q[3] ),
    .S(_05006_),
    .X(_05010_));
 sky130_fd_sc_hd__clkbuf_1 _10353_ (.A(_05010_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _10354_ (.A0(_04730_),
    .A1(\u_rf.reg13_q[4] ),
    .S(_05006_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_1 _10355_ (.A(_05011_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _10356_ (.A0(_04732_),
    .A1(\u_rf.reg13_q[5] ),
    .S(_05006_),
    .X(_05012_));
 sky130_fd_sc_hd__clkbuf_1 _10357_ (.A(_05012_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _10358_ (.A0(_04734_),
    .A1(\u_rf.reg13_q[6] ),
    .S(_05006_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_1 _10359_ (.A(_05013_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _10360_ (.A0(_04736_),
    .A1(\u_rf.reg13_q[7] ),
    .S(_05006_),
    .X(_05014_));
 sky130_fd_sc_hd__clkbuf_1 _10361_ (.A(_05014_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _10362_ (.A0(_04738_),
    .A1(\u_rf.reg13_q[8] ),
    .S(_05006_),
    .X(_05015_));
 sky130_fd_sc_hd__clkbuf_1 _10363_ (.A(_05015_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _10364_ (.A0(_04740_),
    .A1(\u_rf.reg13_q[9] ),
    .S(_05006_),
    .X(_05016_));
 sky130_fd_sc_hd__clkbuf_1 _10365_ (.A(_05016_),
    .X(_00425_));
 sky130_fd_sc_hd__buf_6 _10366_ (.A(_05005_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(_04742_),
    .A1(\u_rf.reg13_q[10] ),
    .S(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__clkbuf_1 _10368_ (.A(_05018_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(_04745_),
    .A1(\u_rf.reg13_q[11] ),
    .S(_05017_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_05019_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(_04747_),
    .A1(\u_rf.reg13_q[12] ),
    .S(_05017_),
    .X(_05020_));
 sky130_fd_sc_hd__clkbuf_1 _10372_ (.A(_05020_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(_04749_),
    .A1(\u_rf.reg13_q[13] ),
    .S(_05017_),
    .X(_05021_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_05021_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(_04751_),
    .A1(\u_rf.reg13_q[14] ),
    .S(_05017_),
    .X(_05022_));
 sky130_fd_sc_hd__clkbuf_1 _10376_ (.A(_05022_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _10377_ (.A0(_04753_),
    .A1(\u_rf.reg13_q[15] ),
    .S(_05017_),
    .X(_05023_));
 sky130_fd_sc_hd__clkbuf_1 _10378_ (.A(_05023_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _10379_ (.A0(_04755_),
    .A1(\u_rf.reg13_q[16] ),
    .S(_05017_),
    .X(_05024_));
 sky130_fd_sc_hd__clkbuf_1 _10380_ (.A(_05024_),
    .X(_00432_));
 sky130_fd_sc_hd__mux2_1 _10381_ (.A0(_04757_),
    .A1(\u_rf.reg13_q[17] ),
    .S(_05017_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(_05025_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(_04759_),
    .A1(\u_rf.reg13_q[18] ),
    .S(_05017_),
    .X(_05026_));
 sky130_fd_sc_hd__clkbuf_1 _10384_ (.A(_05026_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _10385_ (.A0(_04761_),
    .A1(\u_rf.reg13_q[19] ),
    .S(_05017_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_1 _10386_ (.A(_05027_),
    .X(_00435_));
 sky130_fd_sc_hd__clkbuf_8 _10387_ (.A(_05005_),
    .X(_05028_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(_04763_),
    .A1(\u_rf.reg13_q[20] ),
    .S(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_05029_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(_04766_),
    .A1(\u_rf.reg13_q[21] ),
    .S(_05028_),
    .X(_05030_));
 sky130_fd_sc_hd__clkbuf_1 _10391_ (.A(_05030_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(_04768_),
    .A1(\u_rf.reg13_q[22] ),
    .S(_05028_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _10393_ (.A(_05031_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(_04770_),
    .A1(\u_rf.reg13_q[23] ),
    .S(_05028_),
    .X(_05032_));
 sky130_fd_sc_hd__clkbuf_1 _10395_ (.A(_05032_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _10396_ (.A0(_04772_),
    .A1(\u_rf.reg13_q[24] ),
    .S(_05028_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _10397_ (.A(_05033_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _10398_ (.A0(_04774_),
    .A1(\u_rf.reg13_q[25] ),
    .S(_05028_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _10399_ (.A(_05034_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _10400_ (.A0(_04776_),
    .A1(\u_rf.reg13_q[26] ),
    .S(_05028_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_1 _10401_ (.A(_05035_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(_04778_),
    .A1(\u_rf.reg13_q[27] ),
    .S(_05028_),
    .X(_05036_));
 sky130_fd_sc_hd__clkbuf_1 _10403_ (.A(_05036_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(_04780_),
    .A1(\u_rf.reg13_q[28] ),
    .S(_05028_),
    .X(_05037_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_05037_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(_04782_),
    .A1(\u_rf.reg13_q[29] ),
    .S(_05028_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _10407_ (.A(_05038_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(_04784_),
    .A1(\u_rf.reg13_q[30] ),
    .S(_05005_),
    .X(_05039_));
 sky130_fd_sc_hd__clkbuf_1 _10409_ (.A(_05039_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(_04786_),
    .A1(\u_rf.reg13_q[31] ),
    .S(_05005_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_1 _10411_ (.A(_05040_),
    .X(_00447_));
 sky130_fd_sc_hd__or3_4 _10412_ (.A(_04423_),
    .B(_04425_),
    .C(_04936_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_8 _10413_ (.A(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(_04719_),
    .A1(\u_rf.reg14_q[0] ),
    .S(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_05043_),
    .X(_00448_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(_04724_),
    .A1(\u_rf.reg14_q[1] ),
    .S(_05042_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_05044_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(_04726_),
    .A1(\u_rf.reg14_q[2] ),
    .S(_05042_),
    .X(_05045_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_05045_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _10420_ (.A0(_04728_),
    .A1(\u_rf.reg14_q[3] ),
    .S(_05042_),
    .X(_05046_));
 sky130_fd_sc_hd__clkbuf_1 _10421_ (.A(_05046_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(_04730_),
    .A1(\u_rf.reg14_q[4] ),
    .S(_05042_),
    .X(_05047_));
 sky130_fd_sc_hd__clkbuf_1 _10423_ (.A(_05047_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _10424_ (.A0(_04732_),
    .A1(\u_rf.reg14_q[5] ),
    .S(_05042_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_1 _10425_ (.A(_05048_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _10426_ (.A0(_04734_),
    .A1(\u_rf.reg14_q[6] ),
    .S(_05042_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_1 _10427_ (.A(_05049_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _10428_ (.A0(_04736_),
    .A1(\u_rf.reg14_q[7] ),
    .S(_05042_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _10429_ (.A(_05050_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(_04738_),
    .A1(\u_rf.reg14_q[8] ),
    .S(_05042_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _10431_ (.A(_05051_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _10432_ (.A0(_04740_),
    .A1(\u_rf.reg14_q[9] ),
    .S(_05042_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _10433_ (.A(_05052_),
    .X(_00457_));
 sky130_fd_sc_hd__buf_6 _10434_ (.A(_05041_),
    .X(_05053_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(_04742_),
    .A1(\u_rf.reg14_q[10] ),
    .S(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__clkbuf_1 _10436_ (.A(_05054_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(_04745_),
    .A1(\u_rf.reg14_q[11] ),
    .S(_05053_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_05055_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(_04747_),
    .A1(\u_rf.reg14_q[12] ),
    .S(_05053_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_05056_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(_04749_),
    .A1(\u_rf.reg14_q[13] ),
    .S(_05053_),
    .X(_05057_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_05057_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(_04751_),
    .A1(\u_rf.reg14_q[14] ),
    .S(_05053_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_1 _10444_ (.A(_05058_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(_04753_),
    .A1(\u_rf.reg14_q[15] ),
    .S(_05053_),
    .X(_05059_));
 sky130_fd_sc_hd__clkbuf_1 _10446_ (.A(_05059_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(_04755_),
    .A1(\u_rf.reg14_q[16] ),
    .S(_05053_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_1 _10448_ (.A(_05060_),
    .X(_00464_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(_04757_),
    .A1(\u_rf.reg14_q[17] ),
    .S(_05053_),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _10450_ (.A(_05061_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(_04759_),
    .A1(\u_rf.reg14_q[18] ),
    .S(_05053_),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _10452_ (.A(_05062_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(_04761_),
    .A1(\u_rf.reg14_q[19] ),
    .S(_05053_),
    .X(_05063_));
 sky130_fd_sc_hd__clkbuf_1 _10454_ (.A(_05063_),
    .X(_00467_));
 sky130_fd_sc_hd__clkbuf_8 _10455_ (.A(_05041_),
    .X(_05064_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(_04763_),
    .A1(\u_rf.reg14_q[20] ),
    .S(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__clkbuf_1 _10457_ (.A(_05065_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(_04766_),
    .A1(\u_rf.reg14_q[21] ),
    .S(_05064_),
    .X(_05066_));
 sky130_fd_sc_hd__clkbuf_1 _10459_ (.A(_05066_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _10460_ (.A0(_04768_),
    .A1(\u_rf.reg14_q[22] ),
    .S(_05064_),
    .X(_05067_));
 sky130_fd_sc_hd__clkbuf_1 _10461_ (.A(_05067_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(_04770_),
    .A1(\u_rf.reg14_q[23] ),
    .S(_05064_),
    .X(_05068_));
 sky130_fd_sc_hd__clkbuf_1 _10463_ (.A(_05068_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(_04772_),
    .A1(\u_rf.reg14_q[24] ),
    .S(_05064_),
    .X(_05069_));
 sky130_fd_sc_hd__clkbuf_1 _10465_ (.A(_05069_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _10466_ (.A0(_04774_),
    .A1(\u_rf.reg14_q[25] ),
    .S(_05064_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _10467_ (.A(_05070_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _10468_ (.A0(_04776_),
    .A1(\u_rf.reg14_q[26] ),
    .S(_05064_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_1 _10469_ (.A(_05071_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _10470_ (.A0(_04778_),
    .A1(\u_rf.reg14_q[27] ),
    .S(_05064_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_1 _10471_ (.A(_05072_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _10472_ (.A0(_04780_),
    .A1(\u_rf.reg14_q[28] ),
    .S(_05064_),
    .X(_05073_));
 sky130_fd_sc_hd__clkbuf_1 _10473_ (.A(_05073_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _10474_ (.A0(_04782_),
    .A1(\u_rf.reg14_q[29] ),
    .S(_05064_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_1 _10475_ (.A(_05074_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _10476_ (.A0(_04784_),
    .A1(\u_rf.reg14_q[30] ),
    .S(_05041_),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_1 _10477_ (.A(_05075_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _10478_ (.A0(_04786_),
    .A1(\u_rf.reg14_q[31] ),
    .S(_05041_),
    .X(_05076_));
 sky130_fd_sc_hd__clkbuf_1 _10479_ (.A(_05076_),
    .X(_00479_));
 sky130_fd_sc_hd__or3_4 _10480_ (.A(_04423_),
    .B(_04568_),
    .C(_04936_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_8 _10481_ (.A(_05077_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _10482_ (.A0(_04719_),
    .A1(\u_rf.reg15_q[0] ),
    .S(_05078_),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _10483_ (.A(_05079_),
    .X(_00480_));
 sky130_fd_sc_hd__mux2_1 _10484_ (.A0(_04724_),
    .A1(\u_rf.reg15_q[1] ),
    .S(_05078_),
    .X(_05080_));
 sky130_fd_sc_hd__clkbuf_1 _10485_ (.A(_05080_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _10486_ (.A0(_04726_),
    .A1(\u_rf.reg15_q[2] ),
    .S(_05078_),
    .X(_05081_));
 sky130_fd_sc_hd__clkbuf_1 _10487_ (.A(_05081_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _10488_ (.A0(_04728_),
    .A1(\u_rf.reg15_q[3] ),
    .S(_05078_),
    .X(_05082_));
 sky130_fd_sc_hd__clkbuf_1 _10489_ (.A(_05082_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _10490_ (.A0(_04730_),
    .A1(\u_rf.reg15_q[4] ),
    .S(_05078_),
    .X(_05083_));
 sky130_fd_sc_hd__clkbuf_1 _10491_ (.A(_05083_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(_04732_),
    .A1(\u_rf.reg15_q[5] ),
    .S(_05078_),
    .X(_05084_));
 sky130_fd_sc_hd__clkbuf_1 _10493_ (.A(_05084_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(_04734_),
    .A1(\u_rf.reg15_q[6] ),
    .S(_05078_),
    .X(_05085_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_05085_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(_04736_),
    .A1(\u_rf.reg15_q[7] ),
    .S(_05078_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_05086_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(_04738_),
    .A1(\u_rf.reg15_q[8] ),
    .S(_05078_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_05087_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(_04740_),
    .A1(\u_rf.reg15_q[9] ),
    .S(_05078_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_05088_),
    .X(_00489_));
 sky130_fd_sc_hd__buf_6 _10502_ (.A(_05077_),
    .X(_05089_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(_04742_),
    .A1(\u_rf.reg15_q[10] ),
    .S(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _10504_ (.A(_05090_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(_04745_),
    .A1(\u_rf.reg15_q[11] ),
    .S(_05089_),
    .X(_05091_));
 sky130_fd_sc_hd__clkbuf_1 _10506_ (.A(_05091_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(_04747_),
    .A1(\u_rf.reg15_q[12] ),
    .S(_05089_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _10508_ (.A(_05092_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(_04749_),
    .A1(\u_rf.reg15_q[13] ),
    .S(_05089_),
    .X(_05093_));
 sky130_fd_sc_hd__clkbuf_1 _10510_ (.A(_05093_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(_04751_),
    .A1(\u_rf.reg15_q[14] ),
    .S(_05089_),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _10512_ (.A(_05094_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(_04753_),
    .A1(\u_rf.reg15_q[15] ),
    .S(_05089_),
    .X(_05095_));
 sky130_fd_sc_hd__clkbuf_1 _10514_ (.A(_05095_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(_04755_),
    .A1(\u_rf.reg15_q[16] ),
    .S(_05089_),
    .X(_05096_));
 sky130_fd_sc_hd__clkbuf_1 _10516_ (.A(_05096_),
    .X(_00496_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(_04757_),
    .A1(\u_rf.reg15_q[17] ),
    .S(_05089_),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _10518_ (.A(_05097_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(_04759_),
    .A1(\u_rf.reg15_q[18] ),
    .S(_05089_),
    .X(_05098_));
 sky130_fd_sc_hd__clkbuf_1 _10520_ (.A(_05098_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(_04761_),
    .A1(\u_rf.reg15_q[19] ),
    .S(_05089_),
    .X(_05099_));
 sky130_fd_sc_hd__clkbuf_1 _10522_ (.A(_05099_),
    .X(_00499_));
 sky130_fd_sc_hd__buf_6 _10523_ (.A(_05077_),
    .X(_05100_));
 sky130_fd_sc_hd__mux2_1 _10524_ (.A0(_04763_),
    .A1(\u_rf.reg15_q[20] ),
    .S(_05100_),
    .X(_05101_));
 sky130_fd_sc_hd__clkbuf_1 _10525_ (.A(_05101_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(_04766_),
    .A1(\u_rf.reg15_q[21] ),
    .S(_05100_),
    .X(_05102_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(_05102_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(_04768_),
    .A1(\u_rf.reg15_q[22] ),
    .S(_05100_),
    .X(_05103_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(_05103_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(_04770_),
    .A1(\u_rf.reg15_q[23] ),
    .S(_05100_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(_05104_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(_04772_),
    .A1(\u_rf.reg15_q[24] ),
    .S(_05100_),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(_05105_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(_04774_),
    .A1(\u_rf.reg15_q[25] ),
    .S(_05100_),
    .X(_05106_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_05106_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(_04776_),
    .A1(\u_rf.reg15_q[26] ),
    .S(_05100_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_1 _10537_ (.A(_05107_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(_04778_),
    .A1(\u_rf.reg15_q[27] ),
    .S(_05100_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _10539_ (.A(_05108_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(_04780_),
    .A1(\u_rf.reg15_q[28] ),
    .S(_05100_),
    .X(_05109_));
 sky130_fd_sc_hd__clkbuf_1 _10541_ (.A(_05109_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(_04782_),
    .A1(\u_rf.reg15_q[29] ),
    .S(_05100_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_1 _10543_ (.A(_05110_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(_04784_),
    .A1(\u_rf.reg15_q[30] ),
    .S(_05077_),
    .X(_05111_));
 sky130_fd_sc_hd__clkbuf_1 _10545_ (.A(_05111_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(_04786_),
    .A1(\u_rf.reg15_q[31] ),
    .S(_05077_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_05112_),
    .X(_00511_));
 sky130_fd_sc_hd__nand2_1 _10548_ (.A(\u_decod.rf_ff_rd_adr_q_i[4] ),
    .B(\u_decod.rf_write_v_q_i ),
    .Y(_05113_));
 sky130_fd_sc_hd__buf_4 _10549_ (.A(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__nor2_2 _10550_ (.A(_04531_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__clkbuf_8 _10551_ (.A(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(\u_rf.reg16_q[0] ),
    .A1(_04935_),
    .S(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__clkbuf_1 _10553_ (.A(_05117_),
    .X(_00512_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(\u_rf.reg16_q[1] ),
    .A1(_04941_),
    .S(_05116_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_1 _10555_ (.A(_05118_),
    .X(_00513_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(\u_rf.reg16_q[2] ),
    .A1(_04943_),
    .S(_05116_),
    .X(_05119_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(_05119_),
    .X(_00514_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(\u_rf.reg16_q[3] ),
    .A1(_04945_),
    .S(_05116_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_1 _10559_ (.A(_05120_),
    .X(_00515_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\u_rf.reg16_q[4] ),
    .A1(_04947_),
    .S(_05116_),
    .X(_05121_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_05121_),
    .X(_00516_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\u_rf.reg16_q[5] ),
    .A1(_04949_),
    .S(_05116_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(_05122_),
    .X(_00517_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\u_rf.reg16_q[6] ),
    .A1(_04951_),
    .S(_05116_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_05123_),
    .X(_00518_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(\u_rf.reg16_q[7] ),
    .A1(_04953_),
    .S(_05116_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_1 _10567_ (.A(_05124_),
    .X(_00519_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(\u_rf.reg16_q[8] ),
    .A1(_04955_),
    .S(_05116_),
    .X(_05125_));
 sky130_fd_sc_hd__clkbuf_1 _10569_ (.A(_05125_),
    .X(_00520_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\u_rf.reg16_q[9] ),
    .A1(_04957_),
    .S(_05116_),
    .X(_05126_));
 sky130_fd_sc_hd__clkbuf_1 _10571_ (.A(_05126_),
    .X(_00521_));
 sky130_fd_sc_hd__buf_6 _10572_ (.A(_05115_),
    .X(_05127_));
 sky130_fd_sc_hd__mux2_1 _10573_ (.A0(\u_rf.reg16_q[10] ),
    .A1(_04959_),
    .S(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _10574_ (.A(_05128_),
    .X(_00522_));
 sky130_fd_sc_hd__mux2_1 _10575_ (.A0(\u_rf.reg16_q[11] ),
    .A1(_04962_),
    .S(_05127_),
    .X(_05129_));
 sky130_fd_sc_hd__clkbuf_1 _10576_ (.A(_05129_),
    .X(_00523_));
 sky130_fd_sc_hd__mux2_1 _10577_ (.A0(\u_rf.reg16_q[12] ),
    .A1(_04964_),
    .S(_05127_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _10578_ (.A(_05130_),
    .X(_00524_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(\u_rf.reg16_q[13] ),
    .A1(_04966_),
    .S(_05127_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_1 _10580_ (.A(_05131_),
    .X(_00525_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(\u_rf.reg16_q[14] ),
    .A1(_04968_),
    .S(_05127_),
    .X(_05132_));
 sky130_fd_sc_hd__clkbuf_1 _10582_ (.A(_05132_),
    .X(_00526_));
 sky130_fd_sc_hd__mux2_1 _10583_ (.A0(\u_rf.reg16_q[15] ),
    .A1(_04970_),
    .S(_05127_),
    .X(_05133_));
 sky130_fd_sc_hd__clkbuf_1 _10584_ (.A(_05133_),
    .X(_00527_));
 sky130_fd_sc_hd__mux2_1 _10585_ (.A0(\u_rf.reg16_q[16] ),
    .A1(_04972_),
    .S(_05127_),
    .X(_05134_));
 sky130_fd_sc_hd__clkbuf_1 _10586_ (.A(_05134_),
    .X(_00528_));
 sky130_fd_sc_hd__mux2_1 _10587_ (.A0(\u_rf.reg16_q[17] ),
    .A1(_04974_),
    .S(_05127_),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_1 _10588_ (.A(_05135_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _10589_ (.A0(\u_rf.reg16_q[18] ),
    .A1(_04976_),
    .S(_05127_),
    .X(_05136_));
 sky130_fd_sc_hd__clkbuf_1 _10590_ (.A(_05136_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _10591_ (.A0(\u_rf.reg16_q[19] ),
    .A1(_04978_),
    .S(_05127_),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_1 _10592_ (.A(_05137_),
    .X(_00531_));
 sky130_fd_sc_hd__clkbuf_8 _10593_ (.A(_05115_),
    .X(_05138_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\u_rf.reg16_q[20] ),
    .A1(_04980_),
    .S(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__clkbuf_1 _10595_ (.A(_05139_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\u_rf.reg16_q[21] ),
    .A1(_04983_),
    .S(_05138_),
    .X(_05140_));
 sky130_fd_sc_hd__clkbuf_1 _10597_ (.A(_05140_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(\u_rf.reg16_q[22] ),
    .A1(_04985_),
    .S(_05138_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _10599_ (.A(_05141_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\u_rf.reg16_q[23] ),
    .A1(_04987_),
    .S(_05138_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _10601_ (.A(_05142_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(\u_rf.reg16_q[24] ),
    .A1(_04989_),
    .S(_05138_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_1 _10603_ (.A(_05143_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(\u_rf.reg16_q[25] ),
    .A1(_04991_),
    .S(_05138_),
    .X(_05144_));
 sky130_fd_sc_hd__clkbuf_1 _10605_ (.A(_05144_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _10606_ (.A0(\u_rf.reg16_q[26] ),
    .A1(_04993_),
    .S(_05138_),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _10607_ (.A(_05145_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _10608_ (.A0(\u_rf.reg16_q[27] ),
    .A1(_04995_),
    .S(_05138_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_1 _10609_ (.A(_05146_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(\u_rf.reg16_q[28] ),
    .A1(_04997_),
    .S(_05138_),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(_05147_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _10612_ (.A0(\u_rf.reg16_q[29] ),
    .A1(_04999_),
    .S(_05138_),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _10613_ (.A(_05148_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _10614_ (.A0(\u_rf.reg16_q[30] ),
    .A1(_05001_),
    .S(_05115_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_1 _10615_ (.A(_05149_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(\u_rf.reg16_q[31] ),
    .A1(_05003_),
    .S(_05115_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _10617_ (.A(_05150_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_4 _10618_ (.A(_04494_),
    .B(_05114_),
    .Y(_05151_));
 sky130_fd_sc_hd__buf_6 _10619_ (.A(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__mux2_1 _10620_ (.A0(\u_rf.reg17_q[0] ),
    .A1(_04935_),
    .S(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__clkbuf_1 _10621_ (.A(_05153_),
    .X(_00544_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(\u_rf.reg17_q[1] ),
    .A1(_04941_),
    .S(_05152_),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_05154_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _10624_ (.A0(\u_rf.reg17_q[2] ),
    .A1(_04943_),
    .S(_05152_),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_1 _10625_ (.A(_05155_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _10626_ (.A0(\u_rf.reg17_q[3] ),
    .A1(_04945_),
    .S(_05152_),
    .X(_05156_));
 sky130_fd_sc_hd__clkbuf_1 _10627_ (.A(_05156_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(\u_rf.reg17_q[4] ),
    .A1(_04947_),
    .S(_05152_),
    .X(_05157_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_05157_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _10630_ (.A0(\u_rf.reg17_q[5] ),
    .A1(_04949_),
    .S(_05152_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _10631_ (.A(_05158_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _10632_ (.A0(\u_rf.reg17_q[6] ),
    .A1(_04951_),
    .S(_05152_),
    .X(_05159_));
 sky130_fd_sc_hd__clkbuf_1 _10633_ (.A(_05159_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(\u_rf.reg17_q[7] ),
    .A1(_04953_),
    .S(_05152_),
    .X(_05160_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_05160_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _10636_ (.A0(\u_rf.reg17_q[8] ),
    .A1(_04955_),
    .S(_05152_),
    .X(_05161_));
 sky130_fd_sc_hd__clkbuf_1 _10637_ (.A(_05161_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _10638_ (.A0(\u_rf.reg17_q[9] ),
    .A1(_04957_),
    .S(_05152_),
    .X(_05162_));
 sky130_fd_sc_hd__clkbuf_1 _10639_ (.A(_05162_),
    .X(_00553_));
 sky130_fd_sc_hd__buf_8 _10640_ (.A(_05151_),
    .X(_05163_));
 sky130_fd_sc_hd__mux2_1 _10641_ (.A0(\u_rf.reg17_q[10] ),
    .A1(_04959_),
    .S(_05163_),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_1 _10642_ (.A(_05164_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _10643_ (.A0(\u_rf.reg17_q[11] ),
    .A1(_04962_),
    .S(_05163_),
    .X(_05165_));
 sky130_fd_sc_hd__clkbuf_1 _10644_ (.A(_05165_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(\u_rf.reg17_q[12] ),
    .A1(_04964_),
    .S(_05163_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _10646_ (.A(_05166_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _10647_ (.A0(\u_rf.reg17_q[13] ),
    .A1(_04966_),
    .S(_05163_),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _10648_ (.A(_05167_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _10649_ (.A0(\u_rf.reg17_q[14] ),
    .A1(_04968_),
    .S(_05163_),
    .X(_05168_));
 sky130_fd_sc_hd__clkbuf_1 _10650_ (.A(_05168_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _10651_ (.A0(\u_rf.reg17_q[15] ),
    .A1(_04970_),
    .S(_05163_),
    .X(_05169_));
 sky130_fd_sc_hd__clkbuf_1 _10652_ (.A(_05169_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _10653_ (.A0(\u_rf.reg17_q[16] ),
    .A1(_04972_),
    .S(_05163_),
    .X(_05170_));
 sky130_fd_sc_hd__clkbuf_1 _10654_ (.A(_05170_),
    .X(_00560_));
 sky130_fd_sc_hd__mux2_1 _10655_ (.A0(\u_rf.reg17_q[17] ),
    .A1(_04974_),
    .S(_05163_),
    .X(_05171_));
 sky130_fd_sc_hd__clkbuf_1 _10656_ (.A(_05171_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _10657_ (.A0(\u_rf.reg17_q[18] ),
    .A1(_04976_),
    .S(_05163_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_1 _10658_ (.A(_05172_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _10659_ (.A0(\u_rf.reg17_q[19] ),
    .A1(_04978_),
    .S(_05163_),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_1 _10660_ (.A(_05173_),
    .X(_00563_));
 sky130_fd_sc_hd__clkbuf_8 _10661_ (.A(_05151_),
    .X(_05174_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(\u_rf.reg17_q[20] ),
    .A1(_04980_),
    .S(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_05175_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(\u_rf.reg17_q[21] ),
    .A1(_04983_),
    .S(_05174_),
    .X(_05176_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_05176_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(\u_rf.reg17_q[22] ),
    .A1(_04985_),
    .S(_05174_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_05177_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(\u_rf.reg17_q[23] ),
    .A1(_04987_),
    .S(_05174_),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_05178_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(\u_rf.reg17_q[24] ),
    .A1(_04989_),
    .S(_05174_),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_05179_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(\u_rf.reg17_q[25] ),
    .A1(_04991_),
    .S(_05174_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_05180_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(\u_rf.reg17_q[26] ),
    .A1(_04993_),
    .S(_05174_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_05181_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _10676_ (.A0(\u_rf.reg17_q[27] ),
    .A1(_04995_),
    .S(_05174_),
    .X(_05182_));
 sky130_fd_sc_hd__clkbuf_1 _10677_ (.A(_05182_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(\u_rf.reg17_q[28] ),
    .A1(_04997_),
    .S(_05174_),
    .X(_05183_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_05183_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(\u_rf.reg17_q[29] ),
    .A1(_04999_),
    .S(_05174_),
    .X(_05184_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_05184_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(\u_rf.reg17_q[30] ),
    .A1(_05001_),
    .S(_05151_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_05185_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(\u_rf.reg17_q[31] ),
    .A1(_05003_),
    .S(_05151_),
    .X(_05186_));
 sky130_fd_sc_hd__clkbuf_1 _10685_ (.A(_05186_),
    .X(_00575_));
 sky130_fd_sc_hd__nor2_4 _10686_ (.A(_04426_),
    .B(_05114_),
    .Y(_05187_));
 sky130_fd_sc_hd__clkbuf_8 _10687_ (.A(_05187_),
    .X(_05188_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(\u_rf.reg18_q[0] ),
    .A1(_04935_),
    .S(_05188_),
    .X(_05189_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_05189_),
    .X(_00576_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(\u_rf.reg18_q[1] ),
    .A1(_04941_),
    .S(_05188_),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_05190_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(\u_rf.reg18_q[2] ),
    .A1(_04943_),
    .S(_05188_),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_05191_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(\u_rf.reg18_q[3] ),
    .A1(_04945_),
    .S(_05188_),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_05192_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(\u_rf.reg18_q[4] ),
    .A1(_04947_),
    .S(_05188_),
    .X(_05193_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(_05193_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(\u_rf.reg18_q[5] ),
    .A1(_04949_),
    .S(_05188_),
    .X(_05194_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(_05194_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(\u_rf.reg18_q[6] ),
    .A1(_04951_),
    .S(_05188_),
    .X(_05195_));
 sky130_fd_sc_hd__clkbuf_1 _10701_ (.A(_05195_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(\u_rf.reg18_q[7] ),
    .A1(_04953_),
    .S(_05188_),
    .X(_05196_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(_05196_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(\u_rf.reg18_q[8] ),
    .A1(_04955_),
    .S(_05188_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(_05197_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(\u_rf.reg18_q[9] ),
    .A1(_04957_),
    .S(_05188_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_05198_),
    .X(_00585_));
 sky130_fd_sc_hd__buf_8 _10708_ (.A(_05187_),
    .X(_05199_));
 sky130_fd_sc_hd__mux2_1 _10709_ (.A0(\u_rf.reg18_q[10] ),
    .A1(_04959_),
    .S(_05199_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_1 _10710_ (.A(_05200_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _10711_ (.A0(\u_rf.reg18_q[11] ),
    .A1(_04962_),
    .S(_05199_),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_1 _10712_ (.A(_05201_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _10713_ (.A0(\u_rf.reg18_q[12] ),
    .A1(_04964_),
    .S(_05199_),
    .X(_05202_));
 sky130_fd_sc_hd__clkbuf_1 _10714_ (.A(_05202_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _10715_ (.A0(\u_rf.reg18_q[13] ),
    .A1(_04966_),
    .S(_05199_),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_1 _10716_ (.A(_05203_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _10717_ (.A0(\u_rf.reg18_q[14] ),
    .A1(_04968_),
    .S(_05199_),
    .X(_05204_));
 sky130_fd_sc_hd__clkbuf_1 _10718_ (.A(_05204_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _10719_ (.A0(\u_rf.reg18_q[15] ),
    .A1(_04970_),
    .S(_05199_),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_1 _10720_ (.A(_05205_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _10721_ (.A0(\u_rf.reg18_q[16] ),
    .A1(_04972_),
    .S(_05199_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _10722_ (.A(_05206_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _10723_ (.A0(\u_rf.reg18_q[17] ),
    .A1(_04974_),
    .S(_05199_),
    .X(_05207_));
 sky130_fd_sc_hd__clkbuf_1 _10724_ (.A(_05207_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _10725_ (.A0(\u_rf.reg18_q[18] ),
    .A1(_04976_),
    .S(_05199_),
    .X(_05208_));
 sky130_fd_sc_hd__clkbuf_1 _10726_ (.A(_05208_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _10727_ (.A0(\u_rf.reg18_q[19] ),
    .A1(_04978_),
    .S(_05199_),
    .X(_05209_));
 sky130_fd_sc_hd__clkbuf_1 _10728_ (.A(_05209_),
    .X(_00595_));
 sky130_fd_sc_hd__clkbuf_8 _10729_ (.A(_05187_),
    .X(_05210_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(\u_rf.reg18_q[20] ),
    .A1(_04980_),
    .S(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__clkbuf_1 _10731_ (.A(_05211_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(\u_rf.reg18_q[21] ),
    .A1(_04983_),
    .S(_05210_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(_05212_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(\u_rf.reg18_q[22] ),
    .A1(_04985_),
    .S(_05210_),
    .X(_05213_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_05213_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(\u_rf.reg18_q[23] ),
    .A1(_04987_),
    .S(_05210_),
    .X(_05214_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_05214_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(\u_rf.reg18_q[24] ),
    .A1(_04989_),
    .S(_05210_),
    .X(_05215_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_05215_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(\u_rf.reg18_q[25] ),
    .A1(_04991_),
    .S(_05210_),
    .X(_05216_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(_05216_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(\u_rf.reg18_q[26] ),
    .A1(_04993_),
    .S(_05210_),
    .X(_05217_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(_05217_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _10744_ (.A0(\u_rf.reg18_q[27] ),
    .A1(_04995_),
    .S(_05210_),
    .X(_05218_));
 sky130_fd_sc_hd__clkbuf_1 _10745_ (.A(_05218_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(\u_rf.reg18_q[28] ),
    .A1(_04997_),
    .S(_05210_),
    .X(_05219_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_05219_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(\u_rf.reg18_q[29] ),
    .A1(_04999_),
    .S(_05210_),
    .X(_05220_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(_05220_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(\u_rf.reg18_q[30] ),
    .A1(_05001_),
    .S(_05187_),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(_05221_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(\u_rf.reg18_q[31] ),
    .A1(_05003_),
    .S(_05187_),
    .X(_05222_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_05222_),
    .X(_00607_));
 sky130_fd_sc_hd__nor2_2 _10754_ (.A(_04569_),
    .B(_05114_),
    .Y(_05223_));
 sky130_fd_sc_hd__clkbuf_8 _10755_ (.A(_05223_),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(\u_rf.reg19_q[0] ),
    .A1(_04935_),
    .S(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_05225_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(\u_rf.reg19_q[1] ),
    .A1(_04941_),
    .S(_05224_),
    .X(_05226_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_05226_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(\u_rf.reg19_q[2] ),
    .A1(_04943_),
    .S(_05224_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_05227_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(\u_rf.reg19_q[3] ),
    .A1(_04945_),
    .S(_05224_),
    .X(_05228_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_05228_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(\u_rf.reg19_q[4] ),
    .A1(_04947_),
    .S(_05224_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_05229_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(\u_rf.reg19_q[5] ),
    .A1(_04949_),
    .S(_05224_),
    .X(_05230_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_05230_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(\u_rf.reg19_q[6] ),
    .A1(_04951_),
    .S(_05224_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_05231_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(\u_rf.reg19_q[7] ),
    .A1(_04953_),
    .S(_05224_),
    .X(_05232_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_05232_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(\u_rf.reg19_q[8] ),
    .A1(_04955_),
    .S(_05224_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(_05233_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(\u_rf.reg19_q[9] ),
    .A1(_04957_),
    .S(_05224_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_05234_),
    .X(_00617_));
 sky130_fd_sc_hd__clkbuf_8 _10776_ (.A(_05223_),
    .X(_05235_));
 sky130_fd_sc_hd__mux2_1 _10777_ (.A0(\u_rf.reg19_q[10] ),
    .A1(_04959_),
    .S(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__clkbuf_1 _10778_ (.A(_05236_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _10779_ (.A0(\u_rf.reg19_q[11] ),
    .A1(_04962_),
    .S(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__clkbuf_1 _10780_ (.A(_05237_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(\u_rf.reg19_q[12] ),
    .A1(_04964_),
    .S(_05235_),
    .X(_05238_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_05238_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(\u_rf.reg19_q[13] ),
    .A1(_04966_),
    .S(_05235_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_05239_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(\u_rf.reg19_q[14] ),
    .A1(_04968_),
    .S(_05235_),
    .X(_05240_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_05240_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(\u_rf.reg19_q[15] ),
    .A1(_04970_),
    .S(_05235_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_05241_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(\u_rf.reg19_q[16] ),
    .A1(_04972_),
    .S(_05235_),
    .X(_05242_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_05242_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(\u_rf.reg19_q[17] ),
    .A1(_04974_),
    .S(_05235_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_05243_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(\u_rf.reg19_q[18] ),
    .A1(_04976_),
    .S(_05235_),
    .X(_05244_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_05244_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(\u_rf.reg19_q[19] ),
    .A1(_04978_),
    .S(_05235_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_05245_),
    .X(_00627_));
 sky130_fd_sc_hd__buf_6 _10797_ (.A(_05223_),
    .X(_05246_));
 sky130_fd_sc_hd__mux2_1 _10798_ (.A0(\u_rf.reg19_q[20] ),
    .A1(_04980_),
    .S(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__clkbuf_1 _10799_ (.A(_05247_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _10800_ (.A0(\u_rf.reg19_q[21] ),
    .A1(_04983_),
    .S(_05246_),
    .X(_05248_));
 sky130_fd_sc_hd__clkbuf_1 _10801_ (.A(_05248_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _10802_ (.A0(\u_rf.reg19_q[22] ),
    .A1(_04985_),
    .S(_05246_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _10803_ (.A(_05249_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _10804_ (.A0(\u_rf.reg19_q[23] ),
    .A1(_04987_),
    .S(_05246_),
    .X(_05250_));
 sky130_fd_sc_hd__clkbuf_1 _10805_ (.A(_05250_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _10806_ (.A0(\u_rf.reg19_q[24] ),
    .A1(_04989_),
    .S(_05246_),
    .X(_05251_));
 sky130_fd_sc_hd__clkbuf_1 _10807_ (.A(_05251_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(\u_rf.reg19_q[25] ),
    .A1(_04991_),
    .S(_05246_),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_1 _10809_ (.A(_05252_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _10810_ (.A0(\u_rf.reg19_q[26] ),
    .A1(_04993_),
    .S(_05246_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _10811_ (.A(_05253_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _10812_ (.A0(\u_rf.reg19_q[27] ),
    .A1(_04995_),
    .S(_05246_),
    .X(_05254_));
 sky130_fd_sc_hd__clkbuf_1 _10813_ (.A(_05254_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _10814_ (.A0(\u_rf.reg19_q[28] ),
    .A1(_04997_),
    .S(_05246_),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_1 _10815_ (.A(_05255_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _10816_ (.A0(\u_rf.reg19_q[29] ),
    .A1(_04999_),
    .S(_05246_),
    .X(_05256_));
 sky130_fd_sc_hd__clkbuf_1 _10817_ (.A(_05256_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _10818_ (.A0(\u_rf.reg19_q[30] ),
    .A1(_05001_),
    .S(_05223_),
    .X(_05257_));
 sky130_fd_sc_hd__clkbuf_1 _10819_ (.A(_05257_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _10820_ (.A0(\u_rf.reg19_q[31] ),
    .A1(_05003_),
    .S(_05223_),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_1 _10821_ (.A(_05258_),
    .X(_00639_));
 sky130_fd_sc_hd__nor2_2 _10822_ (.A(_04606_),
    .B(_05114_),
    .Y(_05259_));
 sky130_fd_sc_hd__clkbuf_8 _10823_ (.A(_05259_),
    .X(_05260_));
 sky130_fd_sc_hd__mux2_1 _10824_ (.A0(\u_rf.reg20_q[0] ),
    .A1(_04935_),
    .S(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _10825_ (.A(_05261_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _10826_ (.A0(\u_rf.reg20_q[1] ),
    .A1(_04941_),
    .S(_05260_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_1 _10827_ (.A(_05262_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _10828_ (.A0(\u_rf.reg20_q[2] ),
    .A1(_04943_),
    .S(_05260_),
    .X(_05263_));
 sky130_fd_sc_hd__clkbuf_1 _10829_ (.A(_05263_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _10830_ (.A0(\u_rf.reg20_q[3] ),
    .A1(_04945_),
    .S(_05260_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _10831_ (.A(_05264_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _10832_ (.A0(\u_rf.reg20_q[4] ),
    .A1(_04947_),
    .S(_05260_),
    .X(_05265_));
 sky130_fd_sc_hd__clkbuf_1 _10833_ (.A(_05265_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _10834_ (.A0(\u_rf.reg20_q[5] ),
    .A1(_04949_),
    .S(_05260_),
    .X(_05266_));
 sky130_fd_sc_hd__clkbuf_1 _10835_ (.A(_05266_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _10836_ (.A0(\u_rf.reg20_q[6] ),
    .A1(_04951_),
    .S(_05260_),
    .X(_05267_));
 sky130_fd_sc_hd__clkbuf_1 _10837_ (.A(_05267_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _10838_ (.A0(\u_rf.reg20_q[7] ),
    .A1(_04953_),
    .S(_05260_),
    .X(_05268_));
 sky130_fd_sc_hd__clkbuf_1 _10839_ (.A(_05268_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _10840_ (.A0(\u_rf.reg20_q[8] ),
    .A1(_04955_),
    .S(_05260_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_1 _10841_ (.A(_05269_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _10842_ (.A0(\u_rf.reg20_q[9] ),
    .A1(_04957_),
    .S(_05260_),
    .X(_05270_));
 sky130_fd_sc_hd__clkbuf_1 _10843_ (.A(_05270_),
    .X(_00649_));
 sky130_fd_sc_hd__buf_6 _10844_ (.A(_05259_),
    .X(_05271_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(\u_rf.reg20_q[10] ),
    .A1(_04959_),
    .S(_05271_),
    .X(_05272_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_05272_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _10847_ (.A0(\u_rf.reg20_q[11] ),
    .A1(_04962_),
    .S(_05271_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _10848_ (.A(_05273_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(\u_rf.reg20_q[12] ),
    .A1(_04964_),
    .S(_05271_),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_05274_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(\u_rf.reg20_q[13] ),
    .A1(_04966_),
    .S(_05271_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_05275_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(\u_rf.reg20_q[14] ),
    .A1(_04968_),
    .S(_05271_),
    .X(_05276_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_05276_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(\u_rf.reg20_q[15] ),
    .A1(_04970_),
    .S(_05271_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_05277_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(\u_rf.reg20_q[16] ),
    .A1(_04972_),
    .S(_05271_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_05278_),
    .X(_00656_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(\u_rf.reg20_q[17] ),
    .A1(_04974_),
    .S(_05271_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_05279_),
    .X(_00657_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(\u_rf.reg20_q[18] ),
    .A1(_04976_),
    .S(_05271_),
    .X(_05280_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_05280_),
    .X(_00658_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(\u_rf.reg20_q[19] ),
    .A1(_04978_),
    .S(_05271_),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_05281_),
    .X(_00659_));
 sky130_fd_sc_hd__clkbuf_8 _10865_ (.A(_05259_),
    .X(_05282_));
 sky130_fd_sc_hd__mux2_1 _10866_ (.A0(\u_rf.reg20_q[20] ),
    .A1(_04980_),
    .S(_05282_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _10867_ (.A(_05283_),
    .X(_00660_));
 sky130_fd_sc_hd__mux2_1 _10868_ (.A0(\u_rf.reg20_q[21] ),
    .A1(_04983_),
    .S(_05282_),
    .X(_05284_));
 sky130_fd_sc_hd__clkbuf_1 _10869_ (.A(_05284_),
    .X(_00661_));
 sky130_fd_sc_hd__mux2_1 _10870_ (.A0(\u_rf.reg20_q[22] ),
    .A1(_04985_),
    .S(_05282_),
    .X(_05285_));
 sky130_fd_sc_hd__clkbuf_1 _10871_ (.A(_05285_),
    .X(_00662_));
 sky130_fd_sc_hd__mux2_1 _10872_ (.A0(\u_rf.reg20_q[23] ),
    .A1(_04987_),
    .S(_05282_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_1 _10873_ (.A(_05286_),
    .X(_00663_));
 sky130_fd_sc_hd__mux2_1 _10874_ (.A0(\u_rf.reg20_q[24] ),
    .A1(_04989_),
    .S(_05282_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_1 _10875_ (.A(_05287_),
    .X(_00664_));
 sky130_fd_sc_hd__mux2_1 _10876_ (.A0(\u_rf.reg20_q[25] ),
    .A1(_04991_),
    .S(_05282_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _10877_ (.A(_05288_),
    .X(_00665_));
 sky130_fd_sc_hd__mux2_1 _10878_ (.A0(\u_rf.reg20_q[26] ),
    .A1(_04993_),
    .S(_05282_),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_1 _10879_ (.A(_05289_),
    .X(_00666_));
 sky130_fd_sc_hd__mux2_1 _10880_ (.A0(\u_rf.reg20_q[27] ),
    .A1(_04995_),
    .S(_05282_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_1 _10881_ (.A(_05290_),
    .X(_00667_));
 sky130_fd_sc_hd__mux2_1 _10882_ (.A0(\u_rf.reg20_q[28] ),
    .A1(_04997_),
    .S(_05282_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_1 _10883_ (.A(_05291_),
    .X(_00668_));
 sky130_fd_sc_hd__mux2_1 _10884_ (.A0(\u_rf.reg20_q[29] ),
    .A1(_04999_),
    .S(_05282_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _10885_ (.A(_05292_),
    .X(_00669_));
 sky130_fd_sc_hd__mux2_1 _10886_ (.A0(\u_rf.reg20_q[30] ),
    .A1(_05001_),
    .S(_05259_),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_1 _10887_ (.A(_05293_),
    .X(_00670_));
 sky130_fd_sc_hd__mux2_1 _10888_ (.A0(\u_rf.reg20_q[31] ),
    .A1(_05003_),
    .S(_05259_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _10889_ (.A(_05294_),
    .X(_00671_));
 sky130_fd_sc_hd__and2_1 _10890_ (.A(\u_decod.rf_ff_rd_adr_q_i[4] ),
    .B(\u_decod.rf_write_v_q_i ),
    .X(_05295_));
 sky130_fd_sc_hd__and3_2 _10891_ (.A(_04644_),
    .B(_04645_),
    .C(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__buf_6 _10892_ (.A(_05296_),
    .X(_05297_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(\u_rf.reg21_q[0] ),
    .A1(_04935_),
    .S(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_05298_),
    .X(_00672_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(\u_rf.reg21_q[1] ),
    .A1(_04941_),
    .S(_05297_),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_05299_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(\u_rf.reg21_q[2] ),
    .A1(_04943_),
    .S(_05297_),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_05300_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(\u_rf.reg21_q[3] ),
    .A1(_04945_),
    .S(_05297_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_05301_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(\u_rf.reg21_q[4] ),
    .A1(_04947_),
    .S(_05297_),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_05302_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(\u_rf.reg21_q[5] ),
    .A1(_04949_),
    .S(_05297_),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_05303_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(\u_rf.reg21_q[6] ),
    .A1(_04951_),
    .S(_05297_),
    .X(_05304_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_05304_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(\u_rf.reg21_q[7] ),
    .A1(_04953_),
    .S(_05297_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_05305_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(\u_rf.reg21_q[8] ),
    .A1(_04955_),
    .S(_05297_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_05306_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(\u_rf.reg21_q[9] ),
    .A1(_04957_),
    .S(_05297_),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_05307_),
    .X(_00681_));
 sky130_fd_sc_hd__buf_6 _10913_ (.A(_05296_),
    .X(_05308_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(\u_rf.reg21_q[10] ),
    .A1(_04959_),
    .S(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _10915_ (.A(_05309_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _10916_ (.A0(\u_rf.reg21_q[11] ),
    .A1(_04962_),
    .S(_05308_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_1 _10917_ (.A(_05310_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _10918_ (.A0(\u_rf.reg21_q[12] ),
    .A1(_04964_),
    .S(_05308_),
    .X(_05311_));
 sky130_fd_sc_hd__clkbuf_1 _10919_ (.A(_05311_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _10920_ (.A0(\u_rf.reg21_q[13] ),
    .A1(_04966_),
    .S(_05308_),
    .X(_05312_));
 sky130_fd_sc_hd__clkbuf_1 _10921_ (.A(_05312_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(\u_rf.reg21_q[14] ),
    .A1(_04968_),
    .S(_05308_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_05313_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(\u_rf.reg21_q[15] ),
    .A1(_04970_),
    .S(_05308_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_1 _10925_ (.A(_05314_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(\u_rf.reg21_q[16] ),
    .A1(_04972_),
    .S(_05308_),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_1 _10927_ (.A(_05315_),
    .X(_00688_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(\u_rf.reg21_q[17] ),
    .A1(_04974_),
    .S(_05308_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_05316_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _10930_ (.A0(\u_rf.reg21_q[18] ),
    .A1(_04976_),
    .S(_05308_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_1 _10931_ (.A(_05317_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _10932_ (.A0(\u_rf.reg21_q[19] ),
    .A1(_04978_),
    .S(_05308_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _10933_ (.A(_05318_),
    .X(_00691_));
 sky130_fd_sc_hd__buf_6 _10934_ (.A(_05296_),
    .X(_05319_));
 sky130_fd_sc_hd__mux2_1 _10935_ (.A0(\u_rf.reg21_q[20] ),
    .A1(_04980_),
    .S(_05319_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _10936_ (.A(_05320_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(\u_rf.reg21_q[21] ),
    .A1(_04983_),
    .S(_05319_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(_05321_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _10939_ (.A0(\u_rf.reg21_q[22] ),
    .A1(_04985_),
    .S(_05319_),
    .X(_05322_));
 sky130_fd_sc_hd__clkbuf_1 _10940_ (.A(_05322_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _10941_ (.A0(\u_rf.reg21_q[23] ),
    .A1(_04987_),
    .S(_05319_),
    .X(_05323_));
 sky130_fd_sc_hd__clkbuf_1 _10942_ (.A(_05323_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(\u_rf.reg21_q[24] ),
    .A1(_04989_),
    .S(_05319_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_05324_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _10945_ (.A0(\u_rf.reg21_q[25] ),
    .A1(_04991_),
    .S(_05319_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _10946_ (.A(_05325_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _10947_ (.A0(\u_rf.reg21_q[26] ),
    .A1(_04993_),
    .S(_05319_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_1 _10948_ (.A(_05326_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(\u_rf.reg21_q[27] ),
    .A1(_04995_),
    .S(_05319_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_05327_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _10951_ (.A0(\u_rf.reg21_q[28] ),
    .A1(_04997_),
    .S(_05319_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_1 _10952_ (.A(_05328_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _10953_ (.A0(\u_rf.reg21_q[29] ),
    .A1(_04999_),
    .S(_05319_),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _10954_ (.A(_05329_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(\u_rf.reg21_q[30] ),
    .A1(_05001_),
    .S(_05296_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _10956_ (.A(_05330_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _10957_ (.A0(\u_rf.reg21_q[31] ),
    .A1(_05003_),
    .S(_05296_),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _10958_ (.A(_05331_),
    .X(_00703_));
 sky130_fd_sc_hd__and3_4 _10959_ (.A(_04682_),
    .B(_04645_),
    .C(_05295_),
    .X(_05332_));
 sky130_fd_sc_hd__clkbuf_8 _10960_ (.A(_05332_),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(\u_rf.reg22_q[0] ),
    .A1(_04935_),
    .S(_05333_),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_1 _10962_ (.A(_05334_),
    .X(_00704_));
 sky130_fd_sc_hd__mux2_1 _10963_ (.A0(\u_rf.reg22_q[1] ),
    .A1(_04941_),
    .S(_05333_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _10964_ (.A(_05335_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _10965_ (.A0(\u_rf.reg22_q[2] ),
    .A1(_04943_),
    .S(_05333_),
    .X(_05336_));
 sky130_fd_sc_hd__clkbuf_1 _10966_ (.A(_05336_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _10967_ (.A0(\u_rf.reg22_q[3] ),
    .A1(_04945_),
    .S(_05333_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _10968_ (.A(_05337_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _10969_ (.A0(\u_rf.reg22_q[4] ),
    .A1(_04947_),
    .S(_05333_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _10970_ (.A(_05338_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _10971_ (.A0(\u_rf.reg22_q[5] ),
    .A1(_04949_),
    .S(_05333_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _10972_ (.A(_05339_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _10973_ (.A0(\u_rf.reg22_q[6] ),
    .A1(_04951_),
    .S(_05333_),
    .X(_05340_));
 sky130_fd_sc_hd__clkbuf_1 _10974_ (.A(_05340_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _10975_ (.A0(\u_rf.reg22_q[7] ),
    .A1(_04953_),
    .S(_05333_),
    .X(_05341_));
 sky130_fd_sc_hd__clkbuf_1 _10976_ (.A(_05341_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _10977_ (.A0(\u_rf.reg22_q[8] ),
    .A1(_04955_),
    .S(_05333_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_1 _10978_ (.A(_05342_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _10979_ (.A0(\u_rf.reg22_q[9] ),
    .A1(_04957_),
    .S(_05333_),
    .X(_05343_));
 sky130_fd_sc_hd__clkbuf_1 _10980_ (.A(_05343_),
    .X(_00713_));
 sky130_fd_sc_hd__buf_6 _10981_ (.A(_05332_),
    .X(_05344_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(\u_rf.reg22_q[10] ),
    .A1(_04959_),
    .S(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_05345_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(\u_rf.reg22_q[11] ),
    .A1(_04962_),
    .S(_05344_),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_05346_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(\u_rf.reg22_q[12] ),
    .A1(_04964_),
    .S(_05344_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(_05347_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(\u_rf.reg22_q[13] ),
    .A1(_04966_),
    .S(_05344_),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(_05348_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(\u_rf.reg22_q[14] ),
    .A1(_04968_),
    .S(_05344_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(_05349_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(\u_rf.reg22_q[15] ),
    .A1(_04970_),
    .S(_05344_),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(_05350_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(\u_rf.reg22_q[16] ),
    .A1(_04972_),
    .S(_05344_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _10995_ (.A(_05351_),
    .X(_00720_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(\u_rf.reg22_q[17] ),
    .A1(_04974_),
    .S(_05344_),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _10997_ (.A(_05352_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(\u_rf.reg22_q[18] ),
    .A1(_04976_),
    .S(_05344_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _10999_ (.A(_05353_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(\u_rf.reg22_q[19] ),
    .A1(_04978_),
    .S(_05344_),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_1 _11001_ (.A(_05354_),
    .X(_00723_));
 sky130_fd_sc_hd__clkbuf_8 _11002_ (.A(_05332_),
    .X(_05355_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(\u_rf.reg22_q[20] ),
    .A1(_04980_),
    .S(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_05356_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(\u_rf.reg22_q[21] ),
    .A1(_04983_),
    .S(_05355_),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_05357_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(\u_rf.reg22_q[22] ),
    .A1(_04985_),
    .S(_05355_),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_05358_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(\u_rf.reg22_q[23] ),
    .A1(_04987_),
    .S(_05355_),
    .X(_05359_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_05359_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(\u_rf.reg22_q[24] ),
    .A1(_04989_),
    .S(_05355_),
    .X(_05360_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(_05360_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(\u_rf.reg22_q[25] ),
    .A1(_04991_),
    .S(_05355_),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(_05361_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(\u_rf.reg22_q[26] ),
    .A1(_04993_),
    .S(_05355_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _11016_ (.A(_05362_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(\u_rf.reg22_q[27] ),
    .A1(_04995_),
    .S(_05355_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(_05363_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(\u_rf.reg22_q[28] ),
    .A1(_04997_),
    .S(_05355_),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _11020_ (.A(_05364_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(\u_rf.reg22_q[29] ),
    .A1(_04999_),
    .S(_05355_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _11022_ (.A(_05365_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(\u_rf.reg22_q[30] ),
    .A1(_05001_),
    .S(_05332_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _11024_ (.A(_05366_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(\u_rf.reg22_q[31] ),
    .A1(_05003_),
    .S(_05332_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _11026_ (.A(_05367_),
    .X(_00735_));
 sky130_fd_sc_hd__or4_4 _11027_ (.A(_01532_),
    .B(_01536_),
    .C(_04568_),
    .D(_05114_),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_8 _11028_ (.A(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(_04719_),
    .A1(\u_rf.reg23_q[0] ),
    .S(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _11030_ (.A(_05370_),
    .X(_00736_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(_04724_),
    .A1(\u_rf.reg23_q[1] ),
    .S(_05369_),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(_05371_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(_04726_),
    .A1(\u_rf.reg23_q[2] ),
    .S(_05369_),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_05372_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _11035_ (.A0(_04728_),
    .A1(\u_rf.reg23_q[3] ),
    .S(_05369_),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _11036_ (.A(_05373_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(_04730_),
    .A1(\u_rf.reg23_q[4] ),
    .S(_05369_),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(_05374_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(_04732_),
    .A1(\u_rf.reg23_q[5] ),
    .S(_05369_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_05375_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(_04734_),
    .A1(\u_rf.reg23_q[6] ),
    .S(_05369_),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_05376_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(_04736_),
    .A1(\u_rf.reg23_q[7] ),
    .S(_05369_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_05377_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(_04738_),
    .A1(\u_rf.reg23_q[8] ),
    .S(_05369_),
    .X(_05378_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_05378_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(_04740_),
    .A1(\u_rf.reg23_q[9] ),
    .S(_05369_),
    .X(_05379_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_05379_),
    .X(_00745_));
 sky130_fd_sc_hd__buf_6 _11049_ (.A(_05368_),
    .X(_05380_));
 sky130_fd_sc_hd__mux2_1 _11050_ (.A0(_04742_),
    .A1(\u_rf.reg23_q[10] ),
    .S(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _11051_ (.A(_05381_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _11052_ (.A0(_04745_),
    .A1(\u_rf.reg23_q[11] ),
    .S(_05380_),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_1 _11053_ (.A(_05382_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _11054_ (.A0(_04747_),
    .A1(\u_rf.reg23_q[12] ),
    .S(_05380_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _11055_ (.A(_05383_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _11056_ (.A0(_04749_),
    .A1(\u_rf.reg23_q[13] ),
    .S(_05380_),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _11057_ (.A(_05384_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _11058_ (.A0(_04751_),
    .A1(\u_rf.reg23_q[14] ),
    .S(_05380_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _11059_ (.A(_05385_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _11060_ (.A0(_04753_),
    .A1(\u_rf.reg23_q[15] ),
    .S(_05380_),
    .X(_05386_));
 sky130_fd_sc_hd__clkbuf_1 _11061_ (.A(_05386_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _11062_ (.A0(_04755_),
    .A1(\u_rf.reg23_q[16] ),
    .S(_05380_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _11063_ (.A(_05387_),
    .X(_00752_));
 sky130_fd_sc_hd__mux2_1 _11064_ (.A0(_04757_),
    .A1(\u_rf.reg23_q[17] ),
    .S(_05380_),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _11065_ (.A(_05388_),
    .X(_00753_));
 sky130_fd_sc_hd__mux2_1 _11066_ (.A0(_04759_),
    .A1(\u_rf.reg23_q[18] ),
    .S(_05380_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _11067_ (.A(_05389_),
    .X(_00754_));
 sky130_fd_sc_hd__mux2_1 _11068_ (.A0(_04761_),
    .A1(\u_rf.reg23_q[19] ),
    .S(_05380_),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_1 _11069_ (.A(_05390_),
    .X(_00755_));
 sky130_fd_sc_hd__clkbuf_8 _11070_ (.A(_05368_),
    .X(_05391_));
 sky130_fd_sc_hd__mux2_1 _11071_ (.A0(_04763_),
    .A1(\u_rf.reg23_q[20] ),
    .S(_05391_),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _11072_ (.A(_05392_),
    .X(_00756_));
 sky130_fd_sc_hd__mux2_1 _11073_ (.A0(_04766_),
    .A1(\u_rf.reg23_q[21] ),
    .S(_05391_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _11074_ (.A(_05393_),
    .X(_00757_));
 sky130_fd_sc_hd__mux2_1 _11075_ (.A0(_04768_),
    .A1(\u_rf.reg23_q[22] ),
    .S(_05391_),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _11076_ (.A(_05394_),
    .X(_00758_));
 sky130_fd_sc_hd__mux2_1 _11077_ (.A0(_04770_),
    .A1(\u_rf.reg23_q[23] ),
    .S(_05391_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _11078_ (.A(_05395_),
    .X(_00759_));
 sky130_fd_sc_hd__mux2_1 _11079_ (.A0(_04772_),
    .A1(\u_rf.reg23_q[24] ),
    .S(_05391_),
    .X(_05396_));
 sky130_fd_sc_hd__clkbuf_1 _11080_ (.A(_05396_),
    .X(_00760_));
 sky130_fd_sc_hd__mux2_1 _11081_ (.A0(_04774_),
    .A1(\u_rf.reg23_q[25] ),
    .S(_05391_),
    .X(_05397_));
 sky130_fd_sc_hd__clkbuf_1 _11082_ (.A(_05397_),
    .X(_00761_));
 sky130_fd_sc_hd__mux2_1 _11083_ (.A0(_04776_),
    .A1(\u_rf.reg23_q[26] ),
    .S(_05391_),
    .X(_05398_));
 sky130_fd_sc_hd__clkbuf_1 _11084_ (.A(_05398_),
    .X(_00762_));
 sky130_fd_sc_hd__mux2_1 _11085_ (.A0(_04778_),
    .A1(\u_rf.reg23_q[27] ),
    .S(_05391_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _11086_ (.A(_05399_),
    .X(_00763_));
 sky130_fd_sc_hd__mux2_1 _11087_ (.A0(_04780_),
    .A1(\u_rf.reg23_q[28] ),
    .S(_05391_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _11088_ (.A(_05400_),
    .X(_00764_));
 sky130_fd_sc_hd__mux2_1 _11089_ (.A0(_04782_),
    .A1(\u_rf.reg23_q[29] ),
    .S(_05391_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _11090_ (.A(_05401_),
    .X(_00765_));
 sky130_fd_sc_hd__mux2_1 _11091_ (.A0(_04784_),
    .A1(\u_rf.reg23_q[30] ),
    .S(_05368_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _11092_ (.A(_05402_),
    .X(_00766_));
 sky130_fd_sc_hd__mux2_1 _11093_ (.A0(_04786_),
    .A1(\u_rf.reg23_q[31] ),
    .S(_05368_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _11094_ (.A(_05403_),
    .X(_00767_));
 sky130_fd_sc_hd__nor2_4 _11095_ (.A(_04788_),
    .B(_05114_),
    .Y(_05404_));
 sky130_fd_sc_hd__buf_6 _11096_ (.A(_05404_),
    .X(_05405_));
 sky130_fd_sc_hd__mux2_1 _11097_ (.A0(\u_rf.reg24_q[0] ),
    .A1(_04935_),
    .S(_05405_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _11098_ (.A(_05406_),
    .X(_00768_));
 sky130_fd_sc_hd__mux2_1 _11099_ (.A0(\u_rf.reg24_q[1] ),
    .A1(_04941_),
    .S(_05405_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _11100_ (.A(_05407_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _11101_ (.A0(\u_rf.reg24_q[2] ),
    .A1(_04943_),
    .S(_05405_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _11102_ (.A(_05408_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _11103_ (.A0(\u_rf.reg24_q[3] ),
    .A1(_04945_),
    .S(_05405_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _11104_ (.A(_05409_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _11105_ (.A0(\u_rf.reg24_q[4] ),
    .A1(_04947_),
    .S(_05405_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _11106_ (.A(_05410_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(\u_rf.reg24_q[5] ),
    .A1(_04949_),
    .S(_05405_),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _11108_ (.A(_05411_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(\u_rf.reg24_q[6] ),
    .A1(_04951_),
    .S(_05405_),
    .X(_05412_));
 sky130_fd_sc_hd__clkbuf_1 _11110_ (.A(_05412_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(\u_rf.reg24_q[7] ),
    .A1(_04953_),
    .S(_05405_),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _11112_ (.A(_05413_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(\u_rf.reg24_q[8] ),
    .A1(_04955_),
    .S(_05405_),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(_05414_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(\u_rf.reg24_q[9] ),
    .A1(_04957_),
    .S(_05405_),
    .X(_05415_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_05415_),
    .X(_00777_));
 sky130_fd_sc_hd__buf_6 _11117_ (.A(_05404_),
    .X(_05416_));
 sky130_fd_sc_hd__mux2_1 _11118_ (.A0(\u_rf.reg24_q[10] ),
    .A1(_04959_),
    .S(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__clkbuf_1 _11119_ (.A(_05417_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _11120_ (.A0(\u_rf.reg24_q[11] ),
    .A1(_04962_),
    .S(_05416_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _11121_ (.A(_05418_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _11122_ (.A0(\u_rf.reg24_q[12] ),
    .A1(_04964_),
    .S(_05416_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _11123_ (.A(_05419_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _11124_ (.A0(\u_rf.reg24_q[13] ),
    .A1(_04966_),
    .S(_05416_),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _11125_ (.A(_05420_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _11126_ (.A0(\u_rf.reg24_q[14] ),
    .A1(_04968_),
    .S(_05416_),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _11127_ (.A(_05421_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _11128_ (.A0(\u_rf.reg24_q[15] ),
    .A1(_04970_),
    .S(_05416_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _11129_ (.A(_05422_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(\u_rf.reg24_q[16] ),
    .A1(_04972_),
    .S(_05416_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _11131_ (.A(_05423_),
    .X(_00784_));
 sky130_fd_sc_hd__mux2_1 _11132_ (.A0(\u_rf.reg24_q[17] ),
    .A1(_04974_),
    .S(_05416_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_1 _11133_ (.A(_05424_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(\u_rf.reg24_q[18] ),
    .A1(_04976_),
    .S(_05416_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _11135_ (.A(_05425_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(\u_rf.reg24_q[19] ),
    .A1(_04978_),
    .S(_05416_),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_1 _11137_ (.A(_05426_),
    .X(_00787_));
 sky130_fd_sc_hd__clkbuf_8 _11138_ (.A(_05404_),
    .X(_05427_));
 sky130_fd_sc_hd__mux2_1 _11139_ (.A0(\u_rf.reg24_q[20] ),
    .A1(_04980_),
    .S(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_1 _11140_ (.A(_05428_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _11141_ (.A0(\u_rf.reg24_q[21] ),
    .A1(_04983_),
    .S(_05427_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _11142_ (.A(_05429_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _11143_ (.A0(\u_rf.reg24_q[22] ),
    .A1(_04985_),
    .S(_05427_),
    .X(_05430_));
 sky130_fd_sc_hd__clkbuf_1 _11144_ (.A(_05430_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(\u_rf.reg24_q[23] ),
    .A1(_04987_),
    .S(_05427_),
    .X(_05431_));
 sky130_fd_sc_hd__clkbuf_1 _11146_ (.A(_05431_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _11147_ (.A0(\u_rf.reg24_q[24] ),
    .A1(_04989_),
    .S(_05427_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _11148_ (.A(_05432_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _11149_ (.A0(\u_rf.reg24_q[25] ),
    .A1(_04991_),
    .S(_05427_),
    .X(_05433_));
 sky130_fd_sc_hd__clkbuf_1 _11150_ (.A(_05433_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(\u_rf.reg24_q[26] ),
    .A1(_04993_),
    .S(_05427_),
    .X(_05434_));
 sky130_fd_sc_hd__clkbuf_1 _11152_ (.A(_05434_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _11153_ (.A0(\u_rf.reg24_q[27] ),
    .A1(_04995_),
    .S(_05427_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _11154_ (.A(_05435_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _11155_ (.A0(\u_rf.reg24_q[28] ),
    .A1(_04997_),
    .S(_05427_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _11156_ (.A(_05436_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(\u_rf.reg24_q[29] ),
    .A1(_04999_),
    .S(_05427_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(_05437_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _11159_ (.A0(\u_rf.reg24_q[30] ),
    .A1(_05001_),
    .S(_05404_),
    .X(_05438_));
 sky130_fd_sc_hd__clkbuf_1 _11160_ (.A(_05438_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _11161_ (.A0(\u_rf.reg24_q[31] ),
    .A1(_05003_),
    .S(_05404_),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_1 _11162_ (.A(_05439_),
    .X(_00799_));
 sky130_fd_sc_hd__and3_2 _11163_ (.A(_04644_),
    .B(_04825_),
    .C(_05295_),
    .X(_05440_));
 sky130_fd_sc_hd__buf_6 _11164_ (.A(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__mux2_1 _11165_ (.A0(\u_rf.reg25_q[0] ),
    .A1(_04935_),
    .S(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _11166_ (.A(_05442_),
    .X(_00800_));
 sky130_fd_sc_hd__mux2_1 _11167_ (.A0(\u_rf.reg25_q[1] ),
    .A1(_04941_),
    .S(_05441_),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_1 _11168_ (.A(_05443_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(\u_rf.reg25_q[2] ),
    .A1(_04943_),
    .S(_05441_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_05444_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _11171_ (.A0(\u_rf.reg25_q[3] ),
    .A1(_04945_),
    .S(_05441_),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_1 _11172_ (.A(_05445_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _11173_ (.A0(\u_rf.reg25_q[4] ),
    .A1(_04947_),
    .S(_05441_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _11174_ (.A(_05446_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(\u_rf.reg25_q[5] ),
    .A1(_04949_),
    .S(_05441_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_05447_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _11177_ (.A0(\u_rf.reg25_q[6] ),
    .A1(_04951_),
    .S(_05441_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_1 _11178_ (.A(_05448_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _11179_ (.A0(\u_rf.reg25_q[7] ),
    .A1(_04953_),
    .S(_05441_),
    .X(_05449_));
 sky130_fd_sc_hd__clkbuf_1 _11180_ (.A(_05449_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(\u_rf.reg25_q[8] ),
    .A1(_04955_),
    .S(_05441_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_05450_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _11183_ (.A0(\u_rf.reg25_q[9] ),
    .A1(_04957_),
    .S(_05441_),
    .X(_05451_));
 sky130_fd_sc_hd__clkbuf_1 _11184_ (.A(_05451_),
    .X(_00809_));
 sky130_fd_sc_hd__buf_6 _11185_ (.A(_05440_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _11186_ (.A0(\u_rf.reg25_q[10] ),
    .A1(_04959_),
    .S(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _11187_ (.A(_05453_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _11188_ (.A0(\u_rf.reg25_q[11] ),
    .A1(_04962_),
    .S(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _11189_ (.A(_05454_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _11190_ (.A0(\u_rf.reg25_q[12] ),
    .A1(_04964_),
    .S(_05452_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_1 _11191_ (.A(_05455_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _11192_ (.A0(\u_rf.reg25_q[13] ),
    .A1(_04966_),
    .S(_05452_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _11193_ (.A(_05456_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _11194_ (.A0(\u_rf.reg25_q[14] ),
    .A1(_04968_),
    .S(_05452_),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _11195_ (.A(_05457_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _11196_ (.A0(\u_rf.reg25_q[15] ),
    .A1(_04970_),
    .S(_05452_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _11197_ (.A(_05458_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _11198_ (.A0(\u_rf.reg25_q[16] ),
    .A1(_04972_),
    .S(_05452_),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_1 _11199_ (.A(_05459_),
    .X(_00816_));
 sky130_fd_sc_hd__mux2_1 _11200_ (.A0(\u_rf.reg25_q[17] ),
    .A1(_04974_),
    .S(_05452_),
    .X(_05460_));
 sky130_fd_sc_hd__clkbuf_1 _11201_ (.A(_05460_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _11202_ (.A0(\u_rf.reg25_q[18] ),
    .A1(_04976_),
    .S(_05452_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _11203_ (.A(_05461_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _11204_ (.A0(\u_rf.reg25_q[19] ),
    .A1(_04978_),
    .S(_05452_),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_1 _11205_ (.A(_05462_),
    .X(_00819_));
 sky130_fd_sc_hd__clkbuf_8 _11206_ (.A(_05440_),
    .X(_05463_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(\u_rf.reg25_q[20] ),
    .A1(_04980_),
    .S(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_05464_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(\u_rf.reg25_q[21] ),
    .A1(_04983_),
    .S(_05463_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_05465_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(\u_rf.reg25_q[22] ),
    .A1(_04985_),
    .S(_05463_),
    .X(_05466_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(_05466_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(\u_rf.reg25_q[23] ),
    .A1(_04987_),
    .S(_05463_),
    .X(_05467_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(_05467_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(\u_rf.reg25_q[24] ),
    .A1(_04989_),
    .S(_05463_),
    .X(_05468_));
 sky130_fd_sc_hd__clkbuf_1 _11216_ (.A(_05468_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(\u_rf.reg25_q[25] ),
    .A1(_04991_),
    .S(_05463_),
    .X(_05469_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_05469_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(\u_rf.reg25_q[26] ),
    .A1(_04993_),
    .S(_05463_),
    .X(_05470_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_05470_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(\u_rf.reg25_q[27] ),
    .A1(_04995_),
    .S(_05463_),
    .X(_05471_));
 sky130_fd_sc_hd__clkbuf_1 _11222_ (.A(_05471_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _11223_ (.A0(\u_rf.reg25_q[28] ),
    .A1(_04997_),
    .S(_05463_),
    .X(_05472_));
 sky130_fd_sc_hd__clkbuf_1 _11224_ (.A(_05472_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _11225_ (.A0(\u_rf.reg25_q[29] ),
    .A1(_04999_),
    .S(_05463_),
    .X(_05473_));
 sky130_fd_sc_hd__clkbuf_1 _11226_ (.A(_05473_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _11227_ (.A0(\u_rf.reg25_q[30] ),
    .A1(_05001_),
    .S(_05440_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _11228_ (.A(_05474_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _11229_ (.A0(\u_rf.reg25_q[31] ),
    .A1(_05003_),
    .S(_05440_),
    .X(_05475_));
 sky130_fd_sc_hd__clkbuf_1 _11230_ (.A(_05475_),
    .X(_00831_));
 sky130_fd_sc_hd__and3_2 _11231_ (.A(_04682_),
    .B(_04825_),
    .C(_05295_),
    .X(_05476_));
 sky130_fd_sc_hd__buf_6 _11232_ (.A(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _11233_ (.A0(\u_rf.reg26_q[0] ),
    .A1(\u_decod.rf_ff_res_data_i[0] ),
    .S(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_1 _11234_ (.A(_05478_),
    .X(_00832_));
 sky130_fd_sc_hd__mux2_1 _11235_ (.A0(\u_rf.reg26_q[1] ),
    .A1(\u_decod.rf_ff_res_data_i[1] ),
    .S(_05477_),
    .X(_05479_));
 sky130_fd_sc_hd__clkbuf_1 _11236_ (.A(_05479_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _11237_ (.A0(\u_rf.reg26_q[2] ),
    .A1(\u_decod.rf_ff_res_data_i[2] ),
    .S(_05477_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _11238_ (.A(_05480_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(\u_rf.reg26_q[3] ),
    .A1(\u_decod.rf_ff_res_data_i[3] ),
    .S(_05477_),
    .X(_05481_));
 sky130_fd_sc_hd__clkbuf_1 _11240_ (.A(_05481_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(\u_rf.reg26_q[4] ),
    .A1(\u_decod.rf_ff_res_data_i[4] ),
    .S(_05477_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _11242_ (.A(_05482_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _11243_ (.A0(\u_rf.reg26_q[5] ),
    .A1(\u_decod.rf_ff_res_data_i[5] ),
    .S(_05477_),
    .X(_05483_));
 sky130_fd_sc_hd__clkbuf_1 _11244_ (.A(_05483_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _11245_ (.A0(\u_rf.reg26_q[6] ),
    .A1(\u_decod.rf_ff_res_data_i[6] ),
    .S(_05477_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _11246_ (.A(_05484_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _11247_ (.A0(\u_rf.reg26_q[7] ),
    .A1(\u_decod.rf_ff_res_data_i[7] ),
    .S(_05477_),
    .X(_05485_));
 sky130_fd_sc_hd__clkbuf_1 _11248_ (.A(_05485_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _11249_ (.A0(\u_rf.reg26_q[8] ),
    .A1(\u_decod.rf_ff_res_data_i[8] ),
    .S(_05477_),
    .X(_05486_));
 sky130_fd_sc_hd__clkbuf_1 _11250_ (.A(_05486_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _11251_ (.A0(\u_rf.reg26_q[9] ),
    .A1(\u_decod.rf_ff_res_data_i[9] ),
    .S(_05477_),
    .X(_05487_));
 sky130_fd_sc_hd__clkbuf_1 _11252_ (.A(_05487_),
    .X(_00841_));
 sky130_fd_sc_hd__clkbuf_8 _11253_ (.A(_05476_),
    .X(_05488_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(\u_rf.reg26_q[10] ),
    .A1(\u_decod.rf_ff_res_data_i[10] ),
    .S(_05488_),
    .X(_05489_));
 sky130_fd_sc_hd__clkbuf_1 _11255_ (.A(_05489_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(\u_rf.reg26_q[11] ),
    .A1(\u_decod.rf_ff_res_data_i[11] ),
    .S(_05488_),
    .X(_05490_));
 sky130_fd_sc_hd__clkbuf_1 _11257_ (.A(_05490_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _11258_ (.A0(\u_rf.reg26_q[12] ),
    .A1(\u_decod.rf_ff_res_data_i[12] ),
    .S(_05488_),
    .X(_05491_));
 sky130_fd_sc_hd__clkbuf_1 _11259_ (.A(_05491_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(\u_rf.reg26_q[13] ),
    .A1(\u_decod.rf_ff_res_data_i[13] ),
    .S(_05488_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _11261_ (.A(_05492_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(\u_rf.reg26_q[14] ),
    .A1(\u_decod.rf_ff_res_data_i[14] ),
    .S(_05488_),
    .X(_05493_));
 sky130_fd_sc_hd__clkbuf_1 _11263_ (.A(_05493_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(\u_rf.reg26_q[15] ),
    .A1(\u_decod.rf_ff_res_data_i[15] ),
    .S(_05488_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _11265_ (.A(_05494_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(\u_rf.reg26_q[16] ),
    .A1(\u_decod.rf_ff_res_data_i[16] ),
    .S(_05488_),
    .X(_05495_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(_05495_),
    .X(_00848_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(\u_rf.reg26_q[17] ),
    .A1(\u_decod.rf_ff_res_data_i[17] ),
    .S(_05488_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(_05496_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(\u_rf.reg26_q[18] ),
    .A1(\u_decod.rf_ff_res_data_i[18] ),
    .S(_05488_),
    .X(_05497_));
 sky130_fd_sc_hd__clkbuf_1 _11271_ (.A(_05497_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(\u_rf.reg26_q[19] ),
    .A1(\u_decod.rf_ff_res_data_i[19] ),
    .S(_05488_),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _11273_ (.A(_05498_),
    .X(_00851_));
 sky130_fd_sc_hd__clkbuf_8 _11274_ (.A(_05476_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _11275_ (.A0(\u_rf.reg26_q[20] ),
    .A1(\u_decod.rf_ff_res_data_i[20] ),
    .S(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _11276_ (.A(_05500_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _11277_ (.A0(\u_rf.reg26_q[21] ),
    .A1(\u_decod.rf_ff_res_data_i[21] ),
    .S(_05499_),
    .X(_05501_));
 sky130_fd_sc_hd__clkbuf_1 _11278_ (.A(_05501_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _11279_ (.A0(\u_rf.reg26_q[22] ),
    .A1(\u_decod.rf_ff_res_data_i[22] ),
    .S(_05499_),
    .X(_05502_));
 sky130_fd_sc_hd__clkbuf_1 _11280_ (.A(_05502_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _11281_ (.A0(\u_rf.reg26_q[23] ),
    .A1(\u_decod.rf_ff_res_data_i[23] ),
    .S(_05499_),
    .X(_05503_));
 sky130_fd_sc_hd__clkbuf_1 _11282_ (.A(_05503_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _11283_ (.A0(\u_rf.reg26_q[24] ),
    .A1(\u_decod.rf_ff_res_data_i[24] ),
    .S(_05499_),
    .X(_05504_));
 sky130_fd_sc_hd__clkbuf_1 _11284_ (.A(_05504_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _11285_ (.A0(\u_rf.reg26_q[25] ),
    .A1(\u_decod.rf_ff_res_data_i[25] ),
    .S(_05499_),
    .X(_05505_));
 sky130_fd_sc_hd__clkbuf_1 _11286_ (.A(_05505_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _11287_ (.A0(\u_rf.reg26_q[26] ),
    .A1(\u_decod.rf_ff_res_data_i[26] ),
    .S(_05499_),
    .X(_05506_));
 sky130_fd_sc_hd__clkbuf_1 _11288_ (.A(_05506_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _11289_ (.A0(\u_rf.reg26_q[27] ),
    .A1(\u_decod.rf_ff_res_data_i[27] ),
    .S(_05499_),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _11290_ (.A(_05507_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _11291_ (.A0(\u_rf.reg26_q[28] ),
    .A1(\u_decod.rf_ff_res_data_i[28] ),
    .S(_05499_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_1 _11292_ (.A(_05508_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _11293_ (.A0(\u_rf.reg26_q[29] ),
    .A1(\u_decod.rf_ff_res_data_i[29] ),
    .S(_05499_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_1 _11294_ (.A(_05509_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(\u_rf.reg26_q[30] ),
    .A1(\u_decod.rf_ff_res_data_i[30] ),
    .S(_05476_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(_05510_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(\u_rf.reg26_q[31] ),
    .A1(\u_decod.rf_ff_res_data_i[31] ),
    .S(_05476_),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _11298_ (.A(_05511_),
    .X(_00863_));
 sky130_fd_sc_hd__or4_4 _11299_ (.A(_01531_),
    .B(_01535_),
    .C(_04568_),
    .D(_05113_),
    .X(_05512_));
 sky130_fd_sc_hd__clkbuf_8 _11300_ (.A(_05512_),
    .X(_05513_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_04719_),
    .A1(\u_rf.reg27_q[0] ),
    .S(_05513_),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_05514_),
    .X(_00864_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(_04724_),
    .A1(\u_rf.reg27_q[1] ),
    .S(_05513_),
    .X(_05515_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(_05515_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(_04726_),
    .A1(\u_rf.reg27_q[2] ),
    .S(_05513_),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_05516_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(_04728_),
    .A1(\u_rf.reg27_q[3] ),
    .S(_05513_),
    .X(_05517_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_05517_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(_04730_),
    .A1(\u_rf.reg27_q[4] ),
    .S(_05513_),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _11310_ (.A(_05518_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(_04732_),
    .A1(\u_rf.reg27_q[5] ),
    .S(_05513_),
    .X(_05519_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_05519_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(_04734_),
    .A1(\u_rf.reg27_q[6] ),
    .S(_05513_),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_05520_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(_04736_),
    .A1(\u_rf.reg27_q[7] ),
    .S(_05513_),
    .X(_05521_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05521_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(_04738_),
    .A1(\u_rf.reg27_q[8] ),
    .S(_05513_),
    .X(_05522_));
 sky130_fd_sc_hd__clkbuf_1 _11318_ (.A(_05522_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(_04740_),
    .A1(\u_rf.reg27_q[9] ),
    .S(_05513_),
    .X(_05523_));
 sky130_fd_sc_hd__clkbuf_1 _11320_ (.A(_05523_),
    .X(_00873_));
 sky130_fd_sc_hd__buf_6 _11321_ (.A(_05512_),
    .X(_05524_));
 sky130_fd_sc_hd__mux2_1 _11322_ (.A0(_04742_),
    .A1(\u_rf.reg27_q[10] ),
    .S(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__clkbuf_1 _11323_ (.A(_05525_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _11324_ (.A0(_04745_),
    .A1(\u_rf.reg27_q[11] ),
    .S(_05524_),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_1 _11325_ (.A(_05526_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _11326_ (.A0(_04747_),
    .A1(\u_rf.reg27_q[12] ),
    .S(_05524_),
    .X(_05527_));
 sky130_fd_sc_hd__clkbuf_1 _11327_ (.A(_05527_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _11328_ (.A0(_04749_),
    .A1(\u_rf.reg27_q[13] ),
    .S(_05524_),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _11329_ (.A(_05528_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(_04751_),
    .A1(\u_rf.reg27_q[14] ),
    .S(_05524_),
    .X(_05529_));
 sky130_fd_sc_hd__clkbuf_1 _11331_ (.A(_05529_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(_04753_),
    .A1(\u_rf.reg27_q[15] ),
    .S(_05524_),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_1 _11333_ (.A(_05530_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(_04755_),
    .A1(\u_rf.reg27_q[16] ),
    .S(_05524_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _11335_ (.A(_05531_),
    .X(_00880_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(_04757_),
    .A1(\u_rf.reg27_q[17] ),
    .S(_05524_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_1 _11337_ (.A(_05532_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(_04759_),
    .A1(\u_rf.reg27_q[18] ),
    .S(_05524_),
    .X(_05533_));
 sky130_fd_sc_hd__clkbuf_1 _11339_ (.A(_05533_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(_04761_),
    .A1(\u_rf.reg27_q[19] ),
    .S(_05524_),
    .X(_05534_));
 sky130_fd_sc_hd__clkbuf_1 _11341_ (.A(_05534_),
    .X(_00883_));
 sky130_fd_sc_hd__buf_6 _11342_ (.A(_05512_),
    .X(_05535_));
 sky130_fd_sc_hd__mux2_1 _11343_ (.A0(_04763_),
    .A1(\u_rf.reg27_q[20] ),
    .S(_05535_),
    .X(_05536_));
 sky130_fd_sc_hd__clkbuf_1 _11344_ (.A(_05536_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _11345_ (.A0(_04766_),
    .A1(\u_rf.reg27_q[21] ),
    .S(_05535_),
    .X(_05537_));
 sky130_fd_sc_hd__clkbuf_1 _11346_ (.A(_05537_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(_04768_),
    .A1(\u_rf.reg27_q[22] ),
    .S(_05535_),
    .X(_05538_));
 sky130_fd_sc_hd__clkbuf_1 _11348_ (.A(_05538_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _11349_ (.A0(_04770_),
    .A1(\u_rf.reg27_q[23] ),
    .S(_05535_),
    .X(_05539_));
 sky130_fd_sc_hd__clkbuf_1 _11350_ (.A(_05539_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _11351_ (.A0(_04772_),
    .A1(\u_rf.reg27_q[24] ),
    .S(_05535_),
    .X(_05540_));
 sky130_fd_sc_hd__clkbuf_1 _11352_ (.A(_05540_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _11353_ (.A0(_04774_),
    .A1(\u_rf.reg27_q[25] ),
    .S(_05535_),
    .X(_05541_));
 sky130_fd_sc_hd__clkbuf_1 _11354_ (.A(_05541_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(_04776_),
    .A1(\u_rf.reg27_q[26] ),
    .S(_05535_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _11356_ (.A(_05542_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _11357_ (.A0(_04778_),
    .A1(\u_rf.reg27_q[27] ),
    .S(_05535_),
    .X(_05543_));
 sky130_fd_sc_hd__clkbuf_1 _11358_ (.A(_05543_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _11359_ (.A0(_04780_),
    .A1(\u_rf.reg27_q[28] ),
    .S(_05535_),
    .X(_05544_));
 sky130_fd_sc_hd__clkbuf_1 _11360_ (.A(_05544_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _11361_ (.A0(_04782_),
    .A1(\u_rf.reg27_q[29] ),
    .S(_05535_),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _11362_ (.A(_05545_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _11363_ (.A0(_04784_),
    .A1(\u_rf.reg27_q[30] ),
    .S(_05512_),
    .X(_05546_));
 sky130_fd_sc_hd__clkbuf_1 _11364_ (.A(_05546_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(_04786_),
    .A1(\u_rf.reg27_q[31] ),
    .S(_05512_),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _11366_ (.A(_05547_),
    .X(_00895_));
 sky130_fd_sc_hd__nor2_4 _11367_ (.A(_04937_),
    .B(_05114_),
    .Y(_05548_));
 sky130_fd_sc_hd__clkbuf_8 _11368_ (.A(_05548_),
    .X(_05549_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(\u_rf.reg28_q[0] ),
    .A1(\u_decod.rf_ff_res_data_i[0] ),
    .S(_05549_),
    .X(_05550_));
 sky130_fd_sc_hd__clkbuf_1 _11370_ (.A(_05550_),
    .X(_00896_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(\u_rf.reg28_q[1] ),
    .A1(\u_decod.rf_ff_res_data_i[1] ),
    .S(_05549_),
    .X(_05551_));
 sky130_fd_sc_hd__clkbuf_1 _11372_ (.A(_05551_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(\u_rf.reg28_q[2] ),
    .A1(\u_decod.rf_ff_res_data_i[2] ),
    .S(_05549_),
    .X(_05552_));
 sky130_fd_sc_hd__clkbuf_1 _11374_ (.A(_05552_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(\u_rf.reg28_q[3] ),
    .A1(\u_decod.rf_ff_res_data_i[3] ),
    .S(_05549_),
    .X(_05553_));
 sky130_fd_sc_hd__clkbuf_1 _11376_ (.A(_05553_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(\u_rf.reg28_q[4] ),
    .A1(\u_decod.rf_ff_res_data_i[4] ),
    .S(_05549_),
    .X(_05554_));
 sky130_fd_sc_hd__clkbuf_1 _11378_ (.A(_05554_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(\u_rf.reg28_q[5] ),
    .A1(\u_decod.rf_ff_res_data_i[5] ),
    .S(_05549_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _11380_ (.A(_05555_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(\u_rf.reg28_q[6] ),
    .A1(\u_decod.rf_ff_res_data_i[6] ),
    .S(_05549_),
    .X(_05556_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(_05556_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(\u_rf.reg28_q[7] ),
    .A1(\u_decod.rf_ff_res_data_i[7] ),
    .S(_05549_),
    .X(_05557_));
 sky130_fd_sc_hd__clkbuf_1 _11384_ (.A(_05557_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(\u_rf.reg28_q[8] ),
    .A1(\u_decod.rf_ff_res_data_i[8] ),
    .S(_05549_),
    .X(_05558_));
 sky130_fd_sc_hd__clkbuf_1 _11386_ (.A(_05558_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(\u_rf.reg28_q[9] ),
    .A1(\u_decod.rf_ff_res_data_i[9] ),
    .S(_05549_),
    .X(_05559_));
 sky130_fd_sc_hd__clkbuf_1 _11388_ (.A(_05559_),
    .X(_00905_));
 sky130_fd_sc_hd__clkbuf_8 _11389_ (.A(_05548_),
    .X(_05560_));
 sky130_fd_sc_hd__mux2_1 _11390_ (.A0(\u_rf.reg28_q[10] ),
    .A1(\u_decod.rf_ff_res_data_i[10] ),
    .S(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _11391_ (.A(_05561_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _11392_ (.A0(\u_rf.reg28_q[11] ),
    .A1(\u_decod.rf_ff_res_data_i[11] ),
    .S(_05560_),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _11393_ (.A(_05562_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _11394_ (.A0(\u_rf.reg28_q[12] ),
    .A1(\u_decod.rf_ff_res_data_i[12] ),
    .S(_05560_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _11395_ (.A(_05563_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _11396_ (.A0(\u_rf.reg28_q[13] ),
    .A1(\u_decod.rf_ff_res_data_i[13] ),
    .S(_05560_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _11397_ (.A(_05564_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _11398_ (.A0(\u_rf.reg28_q[14] ),
    .A1(\u_decod.rf_ff_res_data_i[14] ),
    .S(_05560_),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _11399_ (.A(_05565_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _11400_ (.A0(\u_rf.reg28_q[15] ),
    .A1(\u_decod.rf_ff_res_data_i[15] ),
    .S(_05560_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _11401_ (.A(_05566_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _11402_ (.A0(\u_rf.reg28_q[16] ),
    .A1(\u_decod.rf_ff_res_data_i[16] ),
    .S(_05560_),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _11403_ (.A(_05567_),
    .X(_00912_));
 sky130_fd_sc_hd__mux2_1 _11404_ (.A0(\u_rf.reg28_q[17] ),
    .A1(\u_decod.rf_ff_res_data_i[17] ),
    .S(_05560_),
    .X(_05568_));
 sky130_fd_sc_hd__clkbuf_1 _11405_ (.A(_05568_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _11406_ (.A0(\u_rf.reg28_q[18] ),
    .A1(\u_decod.rf_ff_res_data_i[18] ),
    .S(_05560_),
    .X(_05569_));
 sky130_fd_sc_hd__clkbuf_1 _11407_ (.A(_05569_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _11408_ (.A0(\u_rf.reg28_q[19] ),
    .A1(\u_decod.rf_ff_res_data_i[19] ),
    .S(_05560_),
    .X(_05570_));
 sky130_fd_sc_hd__clkbuf_1 _11409_ (.A(_05570_),
    .X(_00915_));
 sky130_fd_sc_hd__buf_4 _11410_ (.A(_05548_),
    .X(_05571_));
 sky130_fd_sc_hd__mux2_1 _11411_ (.A0(\u_rf.reg28_q[20] ),
    .A1(\u_decod.rf_ff_res_data_i[20] ),
    .S(_05571_),
    .X(_05572_));
 sky130_fd_sc_hd__clkbuf_1 _11412_ (.A(_05572_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _11413_ (.A0(\u_rf.reg28_q[21] ),
    .A1(\u_decod.rf_ff_res_data_i[21] ),
    .S(_05571_),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _11414_ (.A(_05573_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _11415_ (.A0(\u_rf.reg28_q[22] ),
    .A1(\u_decod.rf_ff_res_data_i[22] ),
    .S(_05571_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _11416_ (.A(_05574_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _11417_ (.A0(\u_rf.reg28_q[23] ),
    .A1(\u_decod.rf_ff_res_data_i[23] ),
    .S(_05571_),
    .X(_05575_));
 sky130_fd_sc_hd__clkbuf_1 _11418_ (.A(_05575_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(\u_rf.reg28_q[24] ),
    .A1(\u_decod.rf_ff_res_data_i[24] ),
    .S(_05571_),
    .X(_05576_));
 sky130_fd_sc_hd__clkbuf_1 _11420_ (.A(_05576_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _11421_ (.A0(\u_rf.reg28_q[25] ),
    .A1(\u_decod.rf_ff_res_data_i[25] ),
    .S(_05571_),
    .X(_05577_));
 sky130_fd_sc_hd__clkbuf_1 _11422_ (.A(_05577_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _11423_ (.A0(\u_rf.reg28_q[26] ),
    .A1(\u_decod.rf_ff_res_data_i[26] ),
    .S(_05571_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _11424_ (.A(_05578_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(\u_rf.reg28_q[27] ),
    .A1(\u_decod.rf_ff_res_data_i[27] ),
    .S(_05571_),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _11426_ (.A(_05579_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(\u_rf.reg28_q[28] ),
    .A1(\u_decod.rf_ff_res_data_i[28] ),
    .S(_05571_),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _11428_ (.A(_05580_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _11429_ (.A0(\u_rf.reg28_q[29] ),
    .A1(\u_decod.rf_ff_res_data_i[29] ),
    .S(_05571_),
    .X(_05581_));
 sky130_fd_sc_hd__clkbuf_1 _11430_ (.A(_05581_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _11431_ (.A0(\u_rf.reg28_q[30] ),
    .A1(\u_decod.rf_ff_res_data_i[30] ),
    .S(_05548_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _11432_ (.A(_05582_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(\u_rf.reg28_q[31] ),
    .A1(\u_decod.rf_ff_res_data_i[31] ),
    .S(_05548_),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _11434_ (.A(_05583_),
    .X(_00927_));
 sky130_fd_sc_hd__or4_4 _11435_ (.A(_01534_),
    .B(_04424_),
    .C(_04936_),
    .D(_05113_),
    .X(_05584_));
 sky130_fd_sc_hd__buf_6 _11436_ (.A(_05584_),
    .X(_05585_));
 sky130_fd_sc_hd__mux2_1 _11437_ (.A0(_04719_),
    .A1(\u_rf.reg29_q[0] ),
    .S(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_1 _11438_ (.A(_05586_),
    .X(_00928_));
 sky130_fd_sc_hd__mux2_1 _11439_ (.A0(_04724_),
    .A1(\u_rf.reg29_q[1] ),
    .S(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__clkbuf_1 _11440_ (.A(_05587_),
    .X(_00929_));
 sky130_fd_sc_hd__mux2_1 _11441_ (.A0(_04726_),
    .A1(\u_rf.reg29_q[2] ),
    .S(_05585_),
    .X(_05588_));
 sky130_fd_sc_hd__clkbuf_1 _11442_ (.A(_05588_),
    .X(_00930_));
 sky130_fd_sc_hd__mux2_1 _11443_ (.A0(_04728_),
    .A1(\u_rf.reg29_q[3] ),
    .S(_05585_),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_1 _11444_ (.A(_05589_),
    .X(_00931_));
 sky130_fd_sc_hd__mux2_1 _11445_ (.A0(_04730_),
    .A1(\u_rf.reg29_q[4] ),
    .S(_05585_),
    .X(_05590_));
 sky130_fd_sc_hd__clkbuf_1 _11446_ (.A(_05590_),
    .X(_00932_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(_04732_),
    .A1(\u_rf.reg29_q[5] ),
    .S(_05585_),
    .X(_05591_));
 sky130_fd_sc_hd__clkbuf_1 _11448_ (.A(_05591_),
    .X(_00933_));
 sky130_fd_sc_hd__mux2_1 _11449_ (.A0(_04734_),
    .A1(\u_rf.reg29_q[6] ),
    .S(_05585_),
    .X(_05592_));
 sky130_fd_sc_hd__clkbuf_1 _11450_ (.A(_05592_),
    .X(_00934_));
 sky130_fd_sc_hd__mux2_1 _11451_ (.A0(_04736_),
    .A1(\u_rf.reg29_q[7] ),
    .S(_05585_),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_1 _11452_ (.A(_05593_),
    .X(_00935_));
 sky130_fd_sc_hd__mux2_1 _11453_ (.A0(_04738_),
    .A1(\u_rf.reg29_q[8] ),
    .S(_05585_),
    .X(_05594_));
 sky130_fd_sc_hd__clkbuf_1 _11454_ (.A(_05594_),
    .X(_00936_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(_04740_),
    .A1(\u_rf.reg29_q[9] ),
    .S(_05585_),
    .X(_05595_));
 sky130_fd_sc_hd__clkbuf_1 _11456_ (.A(_05595_),
    .X(_00937_));
 sky130_fd_sc_hd__buf_6 _11457_ (.A(_05584_),
    .X(_05596_));
 sky130_fd_sc_hd__mux2_1 _11458_ (.A0(_04742_),
    .A1(\u_rf.reg29_q[10] ),
    .S(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__clkbuf_1 _11459_ (.A(_05597_),
    .X(_00938_));
 sky130_fd_sc_hd__mux2_1 _11460_ (.A0(_04745_),
    .A1(\u_rf.reg29_q[11] ),
    .S(_05596_),
    .X(_05598_));
 sky130_fd_sc_hd__clkbuf_1 _11461_ (.A(_05598_),
    .X(_00939_));
 sky130_fd_sc_hd__mux2_1 _11462_ (.A0(_04747_),
    .A1(\u_rf.reg29_q[12] ),
    .S(_05596_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _11463_ (.A(_05599_),
    .X(_00940_));
 sky130_fd_sc_hd__mux2_1 _11464_ (.A0(_04749_),
    .A1(\u_rf.reg29_q[13] ),
    .S(_05596_),
    .X(_05600_));
 sky130_fd_sc_hd__clkbuf_1 _11465_ (.A(_05600_),
    .X(_00941_));
 sky130_fd_sc_hd__mux2_1 _11466_ (.A0(_04751_),
    .A1(\u_rf.reg29_q[14] ),
    .S(_05596_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_1 _11467_ (.A(_05601_),
    .X(_00942_));
 sky130_fd_sc_hd__mux2_1 _11468_ (.A0(_04753_),
    .A1(\u_rf.reg29_q[15] ),
    .S(_05596_),
    .X(_05602_));
 sky130_fd_sc_hd__clkbuf_1 _11469_ (.A(_05602_),
    .X(_00943_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(_04755_),
    .A1(\u_rf.reg29_q[16] ),
    .S(_05596_),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_1 _11471_ (.A(_05603_),
    .X(_00944_));
 sky130_fd_sc_hd__mux2_1 _11472_ (.A0(_04757_),
    .A1(\u_rf.reg29_q[17] ),
    .S(_05596_),
    .X(_05604_));
 sky130_fd_sc_hd__clkbuf_1 _11473_ (.A(_05604_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _11474_ (.A0(_04759_),
    .A1(\u_rf.reg29_q[18] ),
    .S(_05596_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_1 _11475_ (.A(_05605_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(_04761_),
    .A1(\u_rf.reg29_q[19] ),
    .S(_05596_),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_1 _11477_ (.A(_05606_),
    .X(_00947_));
 sky130_fd_sc_hd__buf_6 _11478_ (.A(_05584_),
    .X(_05607_));
 sky130_fd_sc_hd__mux2_1 _11479_ (.A0(_04763_),
    .A1(\u_rf.reg29_q[20] ),
    .S(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_1 _11480_ (.A(_05608_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _11481_ (.A0(_04766_),
    .A1(\u_rf.reg29_q[21] ),
    .S(_05607_),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_1 _11482_ (.A(_05609_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _11483_ (.A0(_04768_),
    .A1(\u_rf.reg29_q[22] ),
    .S(_05607_),
    .X(_05610_));
 sky130_fd_sc_hd__clkbuf_1 _11484_ (.A(_05610_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _11485_ (.A0(_04770_),
    .A1(\u_rf.reg29_q[23] ),
    .S(_05607_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _11486_ (.A(_05611_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _11487_ (.A0(_04772_),
    .A1(\u_rf.reg29_q[24] ),
    .S(_05607_),
    .X(_05612_));
 sky130_fd_sc_hd__clkbuf_1 _11488_ (.A(_05612_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _11489_ (.A0(_04774_),
    .A1(\u_rf.reg29_q[25] ),
    .S(_05607_),
    .X(_05613_));
 sky130_fd_sc_hd__clkbuf_1 _11490_ (.A(_05613_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _11491_ (.A0(_04776_),
    .A1(\u_rf.reg29_q[26] ),
    .S(_05607_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _11492_ (.A(_05614_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _11493_ (.A0(_04778_),
    .A1(\u_rf.reg29_q[27] ),
    .S(_05607_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _11494_ (.A(_05615_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _11495_ (.A0(_04780_),
    .A1(\u_rf.reg29_q[28] ),
    .S(_05607_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _11496_ (.A(_05616_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _11497_ (.A0(_04782_),
    .A1(\u_rf.reg29_q[29] ),
    .S(_05607_),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_1 _11498_ (.A(_05617_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _11499_ (.A0(_04784_),
    .A1(\u_rf.reg29_q[30] ),
    .S(_05584_),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _11500_ (.A(_05618_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _11501_ (.A0(_04786_),
    .A1(\u_rf.reg29_q[31] ),
    .S(_05584_),
    .X(_05619_));
 sky130_fd_sc_hd__clkbuf_1 _11502_ (.A(_05619_),
    .X(_00959_));
 sky130_fd_sc_hd__or3_4 _11503_ (.A(_04425_),
    .B(_04936_),
    .C(_05114_),
    .X(_05620_));
 sky130_fd_sc_hd__buf_6 _11504_ (.A(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(_04719_),
    .A1(\u_rf.reg30_q[0] ),
    .S(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__clkbuf_1 _11506_ (.A(_05622_),
    .X(_00960_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(_04724_),
    .A1(\u_rf.reg30_q[1] ),
    .S(_05621_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_1 _11508_ (.A(_05623_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(_04726_),
    .A1(\u_rf.reg30_q[2] ),
    .S(_05621_),
    .X(_05624_));
 sky130_fd_sc_hd__clkbuf_1 _11510_ (.A(_05624_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(_04728_),
    .A1(\u_rf.reg30_q[3] ),
    .S(_05621_),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_05625_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(_04730_),
    .A1(\u_rf.reg30_q[4] ),
    .S(_05621_),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_1 _11514_ (.A(_05626_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(_04732_),
    .A1(\u_rf.reg30_q[5] ),
    .S(_05621_),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_1 _11516_ (.A(_05627_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(_04734_),
    .A1(\u_rf.reg30_q[6] ),
    .S(_05621_),
    .X(_05628_));
 sky130_fd_sc_hd__clkbuf_1 _11518_ (.A(_05628_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(_04736_),
    .A1(\u_rf.reg30_q[7] ),
    .S(_05621_),
    .X(_05629_));
 sky130_fd_sc_hd__clkbuf_1 _11520_ (.A(_05629_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(_04738_),
    .A1(\u_rf.reg30_q[8] ),
    .S(_05621_),
    .X(_05630_));
 sky130_fd_sc_hd__clkbuf_1 _11522_ (.A(_05630_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(_04740_),
    .A1(\u_rf.reg30_q[9] ),
    .S(_05621_),
    .X(_05631_));
 sky130_fd_sc_hd__clkbuf_1 _11524_ (.A(_05631_),
    .X(_00969_));
 sky130_fd_sc_hd__buf_6 _11525_ (.A(_05620_),
    .X(_05632_));
 sky130_fd_sc_hd__mux2_1 _11526_ (.A0(_04742_),
    .A1(\u_rf.reg30_q[10] ),
    .S(_05632_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_1 _11527_ (.A(_05633_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _11528_ (.A0(_04745_),
    .A1(\u_rf.reg30_q[11] ),
    .S(_05632_),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _11529_ (.A(_05634_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _11530_ (.A0(_04747_),
    .A1(\u_rf.reg30_q[12] ),
    .S(_05632_),
    .X(_05635_));
 sky130_fd_sc_hd__clkbuf_1 _11531_ (.A(_05635_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _11532_ (.A0(_04749_),
    .A1(\u_rf.reg30_q[13] ),
    .S(_05632_),
    .X(_05636_));
 sky130_fd_sc_hd__clkbuf_1 _11533_ (.A(_05636_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _11534_ (.A0(_04751_),
    .A1(\u_rf.reg30_q[14] ),
    .S(_05632_),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _11535_ (.A(_05637_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _11536_ (.A0(_04753_),
    .A1(\u_rf.reg30_q[15] ),
    .S(_05632_),
    .X(_05638_));
 sky130_fd_sc_hd__clkbuf_1 _11537_ (.A(_05638_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _11538_ (.A0(_04755_),
    .A1(\u_rf.reg30_q[16] ),
    .S(_05632_),
    .X(_05639_));
 sky130_fd_sc_hd__clkbuf_1 _11539_ (.A(_05639_),
    .X(_00976_));
 sky130_fd_sc_hd__mux2_1 _11540_ (.A0(_04757_),
    .A1(\u_rf.reg30_q[17] ),
    .S(_05632_),
    .X(_05640_));
 sky130_fd_sc_hd__clkbuf_1 _11541_ (.A(_05640_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _11542_ (.A0(_04759_),
    .A1(\u_rf.reg30_q[18] ),
    .S(_05632_),
    .X(_05641_));
 sky130_fd_sc_hd__clkbuf_1 _11543_ (.A(_05641_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _11544_ (.A0(_04761_),
    .A1(\u_rf.reg30_q[19] ),
    .S(_05632_),
    .X(_05642_));
 sky130_fd_sc_hd__clkbuf_1 _11545_ (.A(_05642_),
    .X(_00979_));
 sky130_fd_sc_hd__clkbuf_8 _11546_ (.A(_05620_),
    .X(_05643_));
 sky130_fd_sc_hd__mux2_1 _11547_ (.A0(_04763_),
    .A1(\u_rf.reg30_q[20] ),
    .S(_05643_),
    .X(_05644_));
 sky130_fd_sc_hd__clkbuf_1 _11548_ (.A(_05644_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _11549_ (.A0(_04766_),
    .A1(\u_rf.reg30_q[21] ),
    .S(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__clkbuf_1 _11550_ (.A(_05645_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _11551_ (.A0(_04768_),
    .A1(\u_rf.reg30_q[22] ),
    .S(_05643_),
    .X(_05646_));
 sky130_fd_sc_hd__clkbuf_1 _11552_ (.A(_05646_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _11553_ (.A0(_04770_),
    .A1(\u_rf.reg30_q[23] ),
    .S(_05643_),
    .X(_05647_));
 sky130_fd_sc_hd__clkbuf_1 _11554_ (.A(_05647_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _11555_ (.A0(_04772_),
    .A1(\u_rf.reg30_q[24] ),
    .S(_05643_),
    .X(_05648_));
 sky130_fd_sc_hd__clkbuf_1 _11556_ (.A(_05648_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _11557_ (.A0(_04774_),
    .A1(\u_rf.reg30_q[25] ),
    .S(_05643_),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_1 _11558_ (.A(_05649_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _11559_ (.A0(_04776_),
    .A1(\u_rf.reg30_q[26] ),
    .S(_05643_),
    .X(_05650_));
 sky130_fd_sc_hd__clkbuf_1 _11560_ (.A(_05650_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _11561_ (.A0(_04778_),
    .A1(\u_rf.reg30_q[27] ),
    .S(_05643_),
    .X(_05651_));
 sky130_fd_sc_hd__clkbuf_1 _11562_ (.A(_05651_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(_04780_),
    .A1(\u_rf.reg30_q[28] ),
    .S(_05643_),
    .X(_05652_));
 sky130_fd_sc_hd__clkbuf_1 _11564_ (.A(_05652_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _11565_ (.A0(_04782_),
    .A1(\u_rf.reg30_q[29] ),
    .S(_05643_),
    .X(_05653_));
 sky130_fd_sc_hd__clkbuf_1 _11566_ (.A(_05653_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _11567_ (.A0(_04784_),
    .A1(\u_rf.reg30_q[30] ),
    .S(_05620_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_1 _11568_ (.A(_05654_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _11569_ (.A0(_04786_),
    .A1(\u_rf.reg30_q[31] ),
    .S(_05620_),
    .X(_05655_));
 sky130_fd_sc_hd__clkbuf_1 _11570_ (.A(_05655_),
    .X(_00991_));
 sky130_fd_sc_hd__or3_4 _11571_ (.A(_04568_),
    .B(_04936_),
    .C(_05114_),
    .X(_05656_));
 sky130_fd_sc_hd__clkbuf_8 _11572_ (.A(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _11573_ (.A0(_04719_),
    .A1(\u_rf.reg31_q[0] ),
    .S(_05657_),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _11574_ (.A(_05658_),
    .X(_00992_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(_04724_),
    .A1(\u_rf.reg31_q[1] ),
    .S(_05657_),
    .X(_05659_));
 sky130_fd_sc_hd__clkbuf_1 _11576_ (.A(_05659_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _11577_ (.A0(_04726_),
    .A1(\u_rf.reg31_q[2] ),
    .S(_05657_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _11578_ (.A(_05660_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _11579_ (.A0(_04728_),
    .A1(\u_rf.reg31_q[3] ),
    .S(_05657_),
    .X(_05661_));
 sky130_fd_sc_hd__clkbuf_1 _11580_ (.A(_05661_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(_04730_),
    .A1(\u_rf.reg31_q[4] ),
    .S(_05657_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _11582_ (.A(_05662_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _11583_ (.A0(_04732_),
    .A1(\u_rf.reg31_q[5] ),
    .S(_05657_),
    .X(_05663_));
 sky130_fd_sc_hd__clkbuf_1 _11584_ (.A(_05663_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _11585_ (.A0(_04734_),
    .A1(\u_rf.reg31_q[6] ),
    .S(_05657_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_1 _11586_ (.A(_05664_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _11587_ (.A0(_04736_),
    .A1(\u_rf.reg31_q[7] ),
    .S(_05657_),
    .X(_05665_));
 sky130_fd_sc_hd__clkbuf_1 _11588_ (.A(_05665_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(_04738_),
    .A1(\u_rf.reg31_q[8] ),
    .S(_05657_),
    .X(_05666_));
 sky130_fd_sc_hd__clkbuf_1 _11590_ (.A(_05666_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(_04740_),
    .A1(\u_rf.reg31_q[9] ),
    .S(_05657_),
    .X(_05667_));
 sky130_fd_sc_hd__clkbuf_1 _11592_ (.A(_05667_),
    .X(_01001_));
 sky130_fd_sc_hd__buf_6 _11593_ (.A(_05656_),
    .X(_05668_));
 sky130_fd_sc_hd__mux2_1 _11594_ (.A0(_04742_),
    .A1(\u_rf.reg31_q[10] ),
    .S(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__clkbuf_1 _11595_ (.A(_05669_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _11596_ (.A0(_04745_),
    .A1(\u_rf.reg31_q[11] ),
    .S(_05668_),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_1 _11597_ (.A(_05670_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _11598_ (.A0(_04747_),
    .A1(\u_rf.reg31_q[12] ),
    .S(_05668_),
    .X(_05671_));
 sky130_fd_sc_hd__clkbuf_1 _11599_ (.A(_05671_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _11600_ (.A0(_04749_),
    .A1(\u_rf.reg31_q[13] ),
    .S(_05668_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _11601_ (.A(_05672_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _11602_ (.A0(_04751_),
    .A1(\u_rf.reg31_q[14] ),
    .S(_05668_),
    .X(_05673_));
 sky130_fd_sc_hd__clkbuf_1 _11603_ (.A(_05673_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _11604_ (.A0(_04753_),
    .A1(\u_rf.reg31_q[15] ),
    .S(_05668_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _11605_ (.A(_05674_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _11606_ (.A0(_04755_),
    .A1(\u_rf.reg31_q[16] ),
    .S(_05668_),
    .X(_05675_));
 sky130_fd_sc_hd__clkbuf_1 _11607_ (.A(_05675_),
    .X(_01008_));
 sky130_fd_sc_hd__mux2_1 _11608_ (.A0(_04757_),
    .A1(\u_rf.reg31_q[17] ),
    .S(_05668_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_1 _11609_ (.A(_05676_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(_04759_),
    .A1(\u_rf.reg31_q[18] ),
    .S(_05668_),
    .X(_05677_));
 sky130_fd_sc_hd__clkbuf_1 _11611_ (.A(_05677_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _11612_ (.A0(_04761_),
    .A1(\u_rf.reg31_q[19] ),
    .S(_05668_),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_1 _11613_ (.A(_05678_),
    .X(_01011_));
 sky130_fd_sc_hd__buf_4 _11614_ (.A(_05656_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(_04763_),
    .A1(\u_rf.reg31_q[20] ),
    .S(_05679_),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _11616_ (.A(_05680_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(_04766_),
    .A1(\u_rf.reg31_q[21] ),
    .S(_05679_),
    .X(_05681_));
 sky130_fd_sc_hd__clkbuf_1 _11618_ (.A(_05681_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(_04768_),
    .A1(\u_rf.reg31_q[22] ),
    .S(_05679_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_05682_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _11621_ (.A0(_04770_),
    .A1(\u_rf.reg31_q[23] ),
    .S(_05679_),
    .X(_05683_));
 sky130_fd_sc_hd__clkbuf_1 _11622_ (.A(_05683_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(_04772_),
    .A1(\u_rf.reg31_q[24] ),
    .S(_05679_),
    .X(_05684_));
 sky130_fd_sc_hd__clkbuf_1 _11624_ (.A(_05684_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _11625_ (.A0(_04774_),
    .A1(\u_rf.reg31_q[25] ),
    .S(_05679_),
    .X(_05685_));
 sky130_fd_sc_hd__clkbuf_1 _11626_ (.A(_05685_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(_04776_),
    .A1(\u_rf.reg31_q[26] ),
    .S(_05679_),
    .X(_05686_));
 sky130_fd_sc_hd__clkbuf_1 _11628_ (.A(_05686_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _11629_ (.A0(_04778_),
    .A1(\u_rf.reg31_q[27] ),
    .S(_05679_),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_1 _11630_ (.A(_05687_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(_04780_),
    .A1(\u_rf.reg31_q[28] ),
    .S(_05679_),
    .X(_05688_));
 sky130_fd_sc_hd__clkbuf_1 _11632_ (.A(_05688_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _11633_ (.A0(_04782_),
    .A1(\u_rf.reg31_q[29] ),
    .S(_05679_),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _11634_ (.A(_05689_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _11635_ (.A0(_04784_),
    .A1(\u_rf.reg31_q[30] ),
    .S(_05656_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_1 _11636_ (.A(_05690_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(_04786_),
    .A1(\u_rf.reg31_q[31] ),
    .S(_05656_),
    .X(_05691_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_05691_),
    .X(_01023_));
 sky130_fd_sc_hd__a22o_1 _11639_ (.A1(\u_decod.dec0.instr_i[7] ),
    .A2(_01227_),
    .B1(_01530_),
    .B2(\u_decod.dec0.instr_i[20] ),
    .X(_05692_));
 sky130_fd_sc_hd__buf_2 _11640_ (.A(net344),
    .X(_05693_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(\u_decod.branch_imm_q_o[0] ),
    .A1(_05692_),
    .S(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__clkbuf_1 _11642_ (.A(_05694_),
    .X(_01024_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(\u_decod.branch_imm_q_o[1] ),
    .A1(_01716_),
    .S(_05693_),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_1 _11644_ (.A(_05695_),
    .X(_01025_));
 sky130_fd_sc_hd__clkbuf_4 _11645_ (.A(net355),
    .X(_05696_));
 sky130_fd_sc_hd__mux2_1 _11646_ (.A0(\u_decod.branch_imm_q_o[2] ),
    .A1(_01774_),
    .S(_05696_),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_1 _11647_ (.A(_05697_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _11648_ (.A0(\u_decod.branch_imm_q_o[3] ),
    .A1(_01831_),
    .S(_05696_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _11649_ (.A(_05698_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _11650_ (.A0(\u_decod.branch_imm_q_o[4] ),
    .A1(_01874_),
    .S(_05696_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _11651_ (.A(_05699_),
    .X(_01028_));
 sky130_fd_sc_hd__buf_2 _11652_ (.A(net345),
    .X(_05700_));
 sky130_fd_sc_hd__and2b_1 _11653_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[5] ),
    .X(_05701_));
 sky130_fd_sc_hd__a31o_1 _11654_ (.A1(\u_decod.dec0.funct7[0] ),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05701_),
    .X(_01029_));
 sky130_fd_sc_hd__and2b_1 _11655_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[6] ),
    .X(_05702_));
 sky130_fd_sc_hd__a31o_1 _11656_ (.A1(\u_decod.dec0.funct7[1] ),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05702_),
    .X(_01030_));
 sky130_fd_sc_hd__and2b_1 _11657_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[7] ),
    .X(_05703_));
 sky130_fd_sc_hd__a31o_1 _11658_ (.A1(\u_decod.dec0.funct7[2] ),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05703_),
    .X(_01031_));
 sky130_fd_sc_hd__and2b_1 _11659_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[8] ),
    .X(_05704_));
 sky130_fd_sc_hd__a31o_1 _11660_ (.A1(\u_decod.dec0.funct7[3] ),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05704_),
    .X(_01032_));
 sky130_fd_sc_hd__and2b_1 _11661_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[9] ),
    .X(_05705_));
 sky130_fd_sc_hd__a31o_1 _11662_ (.A1(\u_decod.dec0.funct7[4] ),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05705_),
    .X(_01033_));
 sky130_fd_sc_hd__and2b_1 _11663_ (.A_N(_05693_),
    .B(\u_decod.branch_imm_q_o[10] ),
    .X(_05706_));
 sky130_fd_sc_hd__a31o_1 _11664_ (.A1(_01079_),
    .A2(_05700_),
    .A3(_02644_),
    .B1(_05706_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _11665_ (.A0(\u_decod.branch_imm_q_o[11] ),
    .A1(_02204_),
    .S(_05696_),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_1 _11666_ (.A(_05707_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _11667_ (.A0(\u_decod.branch_imm_q_o[12] ),
    .A1(_02257_),
    .S(_05696_),
    .X(_05708_));
 sky130_fd_sc_hd__clkbuf_1 _11668_ (.A(_05708_),
    .X(_01036_));
 sky130_fd_sc_hd__nor2_1 _11669_ (.A(_05700_),
    .B(\u_decod.branch_imm_q_o[13] ),
    .Y(_05709_));
 sky130_fd_sc_hd__a21oi_1 _11670_ (.A1(_05700_),
    .A2(_02306_),
    .B1(_05709_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_1 _11671_ (.A(_05693_),
    .B(\u_decod.branch_imm_q_o[14] ),
    .Y(_05710_));
 sky130_fd_sc_hd__a21oi_1 _11672_ (.A1(_05700_),
    .A2(_02391_),
    .B1(_05710_),
    .Y(_01038_));
 sky130_fd_sc_hd__nor2_1 _11673_ (.A(_05693_),
    .B(\u_decod.branch_imm_q_o[15] ),
    .Y(_05711_));
 sky130_fd_sc_hd__a21oi_1 _11674_ (.A1(_05700_),
    .A2(_02418_),
    .B1(_05711_),
    .Y(_01039_));
 sky130_fd_sc_hd__mux2_1 _11675_ (.A0(\u_decod.branch_imm_q_o[16] ),
    .A1(_02465_),
    .S(_05696_),
    .X(_05712_));
 sky130_fd_sc_hd__clkbuf_1 _11676_ (.A(_05712_),
    .X(_01040_));
 sky130_fd_sc_hd__mux2_1 _11677_ (.A0(\u_decod.branch_imm_q_o[17] ),
    .A1(_02509_),
    .S(_05696_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _11678_ (.A(_05713_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _11679_ (.A0(\u_decod.branch_imm_q_o[18] ),
    .A1(_02551_),
    .S(_05696_),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_1 _11680_ (.A(_05714_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _11681_ (.A0(\u_decod.branch_imm_q_o[19] ),
    .A1(_02594_),
    .S(_05696_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _11682_ (.A(_05715_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(\u_decod.branch_imm_q_o[20] ),
    .A1(_02647_),
    .S(_05696_),
    .X(_05716_));
 sky130_fd_sc_hd__clkbuf_1 _11684_ (.A(_05716_),
    .X(_01044_));
 sky130_fd_sc_hd__clkbuf_4 _11685_ (.A(net357),
    .X(_05717_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(\u_decod.branch_imm_q_o[21] ),
    .A1(_02696_),
    .S(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__clkbuf_1 _11687_ (.A(_05718_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(\u_decod.branch_imm_q_o[22] ),
    .A1(_02744_),
    .S(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _11689_ (.A(_05719_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _11690_ (.A0(\u_decod.branch_imm_q_o[23] ),
    .A1(_02792_),
    .S(_05717_),
    .X(_05720_));
 sky130_fd_sc_hd__clkbuf_1 _11691_ (.A(_05720_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(\u_decod.branch_imm_q_o[24] ),
    .A1(_02841_),
    .S(_05717_),
    .X(_05721_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_05721_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(\u_decod.branch_imm_q_o[25] ),
    .A1(_02884_),
    .S(_05717_),
    .X(_05722_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_05722_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(\u_decod.branch_imm_q_o[26] ),
    .A1(_02930_),
    .S(_05717_),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_05723_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(\u_decod.branch_imm_q_o[27] ),
    .A1(_02973_),
    .S(_05717_),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_05724_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(\u_decod.branch_imm_q_o[28] ),
    .A1(_03020_),
    .S(_05717_),
    .X(_05725_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_05725_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(\u_decod.branch_imm_q_o[29] ),
    .A1(_03060_),
    .S(_05717_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_05726_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(\u_decod.branch_imm_q_o[30] ),
    .A1(_03105_),
    .S(_05717_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _11705_ (.A(_05727_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(\u_decod.branch_imm_q_o[31] ),
    .A1(_03143_),
    .S(net346),
    .X(_05728_));
 sky130_fd_sc_hd__clkbuf_1 _11707_ (.A(_05728_),
    .X(_01055_));
 sky130_fd_sc_hd__dfrtp_1 _11708_ (.CLK(clk),
    .D(_00000_),
    .RESET_B(net221),
    .Q(\u_rf.reg2_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11709_ (.CLK(clk),
    .D(_00001_),
    .RESET_B(net236),
    .Q(\u_rf.reg2_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11710_ (.CLK(clk),
    .D(_00002_),
    .RESET_B(net245),
    .Q(\u_rf.reg2_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11711_ (.CLK(clk),
    .D(_00003_),
    .RESET_B(net241),
    .Q(\u_rf.reg2_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11712_ (.CLK(clk),
    .D(_00004_),
    .RESET_B(net227),
    .Q(\u_rf.reg2_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11713_ (.CLK(clk),
    .D(_00005_),
    .RESET_B(net247),
    .Q(\u_rf.reg2_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11714_ (.CLK(clk),
    .D(_00006_),
    .RESET_B(net250),
    .Q(\u_rf.reg2_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11715_ (.CLK(clk),
    .D(_00007_),
    .RESET_B(net234),
    .Q(\u_rf.reg2_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11716_ (.CLK(clk),
    .D(_00008_),
    .RESET_B(net314),
    .Q(\u_rf.reg2_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11717_ (.CLK(clk),
    .D(_00009_),
    .RESET_B(net317),
    .Q(\u_rf.reg2_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11718_ (.CLK(clk),
    .D(_00010_),
    .RESET_B(net247),
    .Q(\u_rf.reg2_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11719_ (.CLK(clk),
    .D(_00011_),
    .RESET_B(net202),
    .Q(\u_rf.reg2_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11720_ (.CLK(clk),
    .D(_00012_),
    .RESET_B(net211),
    .Q(\u_rf.reg2_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11721_ (.CLK(clk),
    .D(_00013_),
    .RESET_B(net281),
    .Q(\u_rf.reg2_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11722_ (.CLK(clk),
    .D(_00014_),
    .RESET_B(net265),
    .Q(\u_rf.reg2_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11723_ (.CLK(clk),
    .D(_00015_),
    .RESET_B(net257),
    .Q(\u_rf.reg2_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11724_ (.CLK(clk),
    .D(_00016_),
    .RESET_B(net223),
    .Q(\u_rf.reg2_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11725_ (.CLK(clk),
    .D(_00017_),
    .RESET_B(net280),
    .Q(\u_rf.reg2_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11726_ (.CLK(clk),
    .D(_00018_),
    .RESET_B(net215),
    .Q(\u_rf.reg2_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11727_ (.CLK(clk),
    .D(_00019_),
    .RESET_B(net216),
    .Q(\u_rf.reg2_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11728_ (.CLK(clk),
    .D(_00020_),
    .RESET_B(net271),
    .Q(\u_rf.reg2_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11729_ (.CLK(clk),
    .D(_00021_),
    .RESET_B(net271),
    .Q(\u_rf.reg2_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11730_ (.CLK(clk),
    .D(_00022_),
    .RESET_B(net286),
    .Q(\u_rf.reg2_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11731_ (.CLK(clk),
    .D(_00023_),
    .RESET_B(net277),
    .Q(\u_rf.reg2_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11732_ (.CLK(clk),
    .D(_00024_),
    .RESET_B(net349),
    .Q(\u_rf.reg2_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11733_ (.CLK(clk),
    .D(_00025_),
    .RESET_B(net262),
    .Q(\u_rf.reg2_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11734_ (.CLK(clk),
    .D(_00026_),
    .RESET_B(net296),
    .Q(\u_rf.reg2_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11735_ (.CLK(clk),
    .D(_00027_),
    .RESET_B(net307),
    .Q(\u_rf.reg2_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11736_ (.CLK(clk),
    .D(_00028_),
    .RESET_B(net353),
    .Q(\u_rf.reg2_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11737_ (.CLK(clk),
    .D(_00029_),
    .RESET_B(net355),
    .Q(\u_rf.reg2_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11738_ (.CLK(clk),
    .D(_00030_),
    .RESET_B(net343),
    .Q(\u_rf.reg2_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11739_ (.CLK(clk),
    .D(_00031_),
    .RESET_B(net343),
    .Q(\u_rf.reg2_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11740_ (.CLK(clk),
    .D(_00032_),
    .RESET_B(net245),
    .Q(\u_rf.reg1_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11741_ (.CLK(clk),
    .D(_00033_),
    .RESET_B(net236),
    .Q(\u_rf.reg1_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11742_ (.CLK(clk),
    .D(_00034_),
    .RESET_B(net245),
    .Q(\u_rf.reg1_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11743_ (.CLK(clk),
    .D(_00035_),
    .RESET_B(net243),
    .Q(\u_rf.reg1_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11744_ (.CLK(clk),
    .D(_00036_),
    .RESET_B(net227),
    .Q(\u_rf.reg1_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11745_ (.CLK(clk),
    .D(_00037_),
    .RESET_B(net324),
    .Q(\u_rf.reg1_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11746_ (.CLK(clk),
    .D(_00038_),
    .RESET_B(net251),
    .Q(\u_rf.reg1_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11747_ (.CLK(clk),
    .D(_00039_),
    .RESET_B(net234),
    .Q(\u_rf.reg1_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11748_ (.CLK(clk),
    .D(_00040_),
    .RESET_B(net312),
    .Q(\u_rf.reg1_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11749_ (.CLK(clk),
    .D(_00041_),
    .RESET_B(net312),
    .Q(\u_rf.reg1_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11750_ (.CLK(clk),
    .D(_00042_),
    .RESET_B(net247),
    .Q(\u_rf.reg1_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11751_ (.CLK(clk),
    .D(_00043_),
    .RESET_B(net202),
    .Q(\u_rf.reg1_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11752_ (.CLK(clk),
    .D(_00044_),
    .RESET_B(net211),
    .Q(\u_rf.reg1_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11753_ (.CLK(clk),
    .D(_00045_),
    .RESET_B(net288),
    .Q(\u_rf.reg1_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11754_ (.CLK(clk),
    .D(_00046_),
    .RESET_B(net265),
    .Q(\u_rf.reg1_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11755_ (.CLK(clk),
    .D(_00047_),
    .RESET_B(net257),
    .Q(\u_rf.reg1_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11756_ (.CLK(clk),
    .D(_00048_),
    .RESET_B(net221),
    .Q(\u_rf.reg1_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11757_ (.CLK(clk),
    .D(_00049_),
    .RESET_B(net280),
    .Q(\u_rf.reg1_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11758_ (.CLK(clk),
    .D(_00050_),
    .RESET_B(net215),
    .Q(\u_rf.reg1_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11759_ (.CLK(clk),
    .D(_00051_),
    .RESET_B(net256),
    .Q(\u_rf.reg1_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11760_ (.CLK(clk),
    .D(_00052_),
    .RESET_B(net272),
    .Q(\u_rf.reg1_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11761_ (.CLK(clk),
    .D(_00053_),
    .RESET_B(net271),
    .Q(\u_rf.reg1_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11762_ (.CLK(clk),
    .D(_00054_),
    .RESET_B(net291),
    .Q(\u_rf.reg1_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11763_ (.CLK(clk),
    .D(_00055_),
    .RESET_B(net277),
    .Q(\u_rf.reg1_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11764_ (.CLK(clk),
    .D(_00056_),
    .RESET_B(net349),
    .Q(\u_rf.reg1_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11765_ (.CLK(clk),
    .D(_00057_),
    .RESET_B(net263),
    .Q(\u_rf.reg1_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11766_ (.CLK(clk),
    .D(_00058_),
    .RESET_B(net300),
    .Q(\u_rf.reg1_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11767_ (.CLK(clk),
    .D(_00059_),
    .RESET_B(net306),
    .Q(\u_rf.reg1_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11768_ (.CLK(clk),
    .D(_00060_),
    .RESET_B(net358),
    .Q(\u_rf.reg1_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11769_ (.CLK(clk),
    .D(_00061_),
    .RESET_B(net355),
    .Q(\u_rf.reg1_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11770_ (.CLK(clk),
    .D(_00062_),
    .RESET_B(net341),
    .Q(\u_rf.reg1_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11771_ (.CLK(clk),
    .D(_00063_),
    .RESET_B(net339),
    .Q(\u_rf.reg1_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11772_ (.CLK(clk),
    .D(net369),
    .RESET_B(net369),
    .Q(\u_ifetch.reset_n_q ));
 sky130_fd_sc_hd__dfrtp_2 _11773_ (.CLK(clk),
    .D(net134),
    .RESET_B(net360),
    .Q(\u_decod.pc0_q_i[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11774_ (.CLK(clk),
    .D(net145),
    .RESET_B(net360),
    .Q(\u_decod.pc0_q_i[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11775_ (.CLK(clk),
    .D(net156),
    .RESET_B(net360),
    .Q(\u_decod.pc0_q_i[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11776_ (.CLK(clk),
    .D(net159),
    .RESET_B(net361),
    .Q(\u_decod.pc0_q_i[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11777_ (.CLK(clk),
    .D(net160),
    .RESET_B(net362),
    .Q(\u_decod.pc0_q_i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11778_ (.CLK(clk),
    .D(net161),
    .RESET_B(net362),
    .Q(\u_decod.pc0_q_i[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11779_ (.CLK(clk),
    .D(net162),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11780_ (.CLK(clk),
    .D(net163),
    .RESET_B(net363),
    .Q(\u_decod.pc0_q_i[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11781_ (.CLK(clk),
    .D(net164),
    .RESET_B(net363),
    .Q(\u_decod.pc0_q_i[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11782_ (.CLK(clk),
    .D(net165),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11783_ (.CLK(clk),
    .D(net135),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11784_ (.CLK(clk),
    .D(net136),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[11] ));
 sky130_fd_sc_hd__dfrtp_2 _11785_ (.CLK(clk),
    .D(net137),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11786_ (.CLK(clk),
    .D(net138),
    .RESET_B(net364),
    .Q(\u_decod.pc0_q_i[13] ));
 sky130_fd_sc_hd__dfrtp_2 _11787_ (.CLK(clk),
    .D(net139),
    .RESET_B(net365),
    .Q(\u_decod.pc0_q_i[14] ));
 sky130_fd_sc_hd__dfrtp_2 _11788_ (.CLK(clk),
    .D(net140),
    .RESET_B(net365),
    .Q(\u_decod.pc0_q_i[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11789_ (.CLK(clk),
    .D(net141),
    .RESET_B(net365),
    .Q(\u_decod.pc0_q_i[16] ));
 sky130_fd_sc_hd__dfrtp_2 _11790_ (.CLK(clk),
    .D(net142),
    .RESET_B(net365),
    .Q(\u_decod.pc0_q_i[17] ));
 sky130_fd_sc_hd__dfrtp_4 _11791_ (.CLK(clk),
    .D(net143),
    .RESET_B(net371),
    .Q(\u_decod.pc0_q_i[18] ));
 sky130_fd_sc_hd__dfrtp_2 _11792_ (.CLK(clk),
    .D(net144),
    .RESET_B(net371),
    .Q(\u_decod.pc0_q_i[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11793_ (.CLK(clk),
    .D(net146),
    .RESET_B(net371),
    .Q(\u_decod.pc0_q_i[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11794_ (.CLK(clk),
    .D(net147),
    .RESET_B(net370),
    .Q(\u_decod.pc0_q_i[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11795_ (.CLK(clk),
    .D(net148),
    .RESET_B(net370),
    .Q(\u_decod.pc0_q_i[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11796_ (.CLK(clk),
    .D(net149),
    .RESET_B(net370),
    .Q(\u_decod.pc0_q_i[23] ));
 sky130_fd_sc_hd__dfrtp_2 _11797_ (.CLK(clk),
    .D(net150),
    .RESET_B(net372),
    .Q(\u_decod.pc0_q_i[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11798_ (.CLK(clk),
    .D(net151),
    .RESET_B(net370),
    .Q(\u_decod.pc0_q_i[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11799_ (.CLK(clk),
    .D(net152),
    .RESET_B(net369),
    .Q(\u_decod.pc0_q_i[26] ));
 sky130_fd_sc_hd__dfrtp_2 _11800_ (.CLK(clk),
    .D(net153),
    .RESET_B(net369),
    .Q(\u_decod.pc0_q_i[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11801_ (.CLK(clk),
    .D(net154),
    .RESET_B(net368),
    .Q(\u_decod.pc0_q_i[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11802_ (.CLK(clk),
    .D(net155),
    .RESET_B(net368),
    .Q(\u_decod.pc0_q_i[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11803_ (.CLK(clk),
    .D(net157),
    .RESET_B(net368),
    .Q(\u_decod.pc0_q_i[30] ));
 sky130_fd_sc_hd__dfrtp_2 _11804_ (.CLK(clk),
    .D(net158),
    .RESET_B(net361),
    .Q(\u_decod.pc0_q_i[31] ));
 sky130_fd_sc_hd__dfrtp_2 _11805_ (.CLK(clk),
    .D(net1),
    .RESET_B(net320),
    .Q(\u_decod.dec0.instr_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11806_ (.CLK(clk),
    .D(net12),
    .RESET_B(net320),
    .Q(\u_decod.dec0.instr_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11807_ (.CLK(clk),
    .D(net23),
    .RESET_B(net320),
    .Q(\u_decod.dec0.instr_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11808_ (.CLK(clk),
    .D(net26),
    .RESET_B(net320),
    .Q(\u_decod.dec0.instr_i[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11809_ (.CLK(clk),
    .D(net27),
    .RESET_B(net319),
    .Q(\u_decod.dec0.instr_i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11810_ (.CLK(clk),
    .D(net28),
    .RESET_B(net320),
    .Q(\u_decod.dec0.instr_i[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11811_ (.CLK(clk),
    .D(net29),
    .RESET_B(net319),
    .Q(\u_decod.dec0.instr_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11812_ (.CLK(clk),
    .D(net30),
    .RESET_B(net321),
    .Q(\u_decod.dec0.instr_i[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11813_ (.CLK(clk),
    .D(net31),
    .RESET_B(net331),
    .Q(\u_decod.dec0.instr_i[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11814_ (.CLK(clk),
    .D(net32),
    .RESET_B(net331),
    .Q(\u_decod.dec0.instr_i[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11815_ (.CLK(clk),
    .D(net2),
    .RESET_B(net328),
    .Q(\u_decod.dec0.instr_i[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11816_ (.CLK(clk),
    .D(net3),
    .RESET_B(net331),
    .Q(\u_decod.dec0.instr_i[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11817_ (.CLK(clk),
    .D(net4),
    .RESET_B(net319),
    .Q(\u_decod.dec0.funct3[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11818_ (.CLK(clk),
    .D(net5),
    .RESET_B(net319),
    .Q(\u_decod.dec0.funct3[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11819_ (.CLK(clk),
    .D(net6),
    .RESET_B(net319),
    .Q(\u_decod.dec0.funct3[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11820_ (.CLK(clk),
    .D(net7),
    .RESET_B(net339),
    .Q(\u_decod.dec0.instr_i[15] ));
 sky130_fd_sc_hd__dfrtp_4 _11821_ (.CLK(clk),
    .D(net8),
    .RESET_B(net339),
    .Q(\u_decod.dec0.instr_i[16] ));
 sky130_fd_sc_hd__dfrtp_4 _11822_ (.CLK(clk),
    .D(net9),
    .RESET_B(net344),
    .Q(\u_decod.dec0.instr_i[17] ));
 sky130_fd_sc_hd__dfrtp_4 _11823_ (.CLK(clk),
    .D(net10),
    .RESET_B(net344),
    .Q(\u_decod.dec0.instr_i[18] ));
 sky130_fd_sc_hd__dfrtp_4 _11824_ (.CLK(clk),
    .D(net11),
    .RESET_B(net344),
    .Q(\u_decod.dec0.instr_i[19] ));
 sky130_fd_sc_hd__dfrtp_4 _11825_ (.CLK(clk),
    .D(net13),
    .RESET_B(net321),
    .Q(\u_decod.dec0.instr_i[20] ));
 sky130_fd_sc_hd__dfrtp_4 _11826_ (.CLK(clk),
    .D(net14),
    .RESET_B(net328),
    .Q(\u_decod.dec0.instr_i[21] ));
 sky130_fd_sc_hd__dfrtp_4 _11827_ (.CLK(clk),
    .D(net15),
    .RESET_B(net328),
    .Q(\u_decod.dec0.instr_i[22] ));
 sky130_fd_sc_hd__dfrtp_4 _11828_ (.CLK(clk),
    .D(net16),
    .RESET_B(net328),
    .Q(\u_decod.dec0.instr_i[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11829_ (.CLK(clk),
    .D(net17),
    .RESET_B(net323),
    .Q(\u_decod.dec0.instr_i[24] ));
 sky130_fd_sc_hd__dfrtp_2 _11830_ (.CLK(clk),
    .D(net18),
    .RESET_B(net329),
    .Q(\u_decod.dec0.funct7[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11831_ (.CLK(clk),
    .D(net19),
    .RESET_B(net329),
    .Q(\u_decod.dec0.funct7[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11832_ (.CLK(clk),
    .D(net20),
    .RESET_B(net321),
    .Q(\u_decod.dec0.funct7[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11833_ (.CLK(clk),
    .D(net21),
    .RESET_B(net321),
    .Q(\u_decod.dec0.funct7[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11834_ (.CLK(clk),
    .D(net22),
    .RESET_B(net322),
    .Q(\u_decod.dec0.funct7[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11835_ (.CLK(clk),
    .D(net24),
    .RESET_B(net328),
    .Q(\u_decod.dec0.funct7[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11836_ (.CLK(clk),
    .D(net25),
    .RESET_B(net321),
    .Q(\u_decod.dec0.funct7[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11837_ (.CLK(clk),
    .D(_00064_),
    .RESET_B(net244),
    .Q(\u_rf.reg0_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11838_ (.CLK(clk),
    .D(_00065_),
    .RESET_B(net236),
    .Q(\u_rf.reg0_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11839_ (.CLK(clk),
    .D(_00066_),
    .RESET_B(net241),
    .Q(\u_rf.reg0_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11840_ (.CLK(clk),
    .D(_00067_),
    .RESET_B(net231),
    .Q(\u_rf.reg0_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11841_ (.CLK(clk),
    .D(_00068_),
    .RESET_B(net227),
    .Q(\u_rf.reg0_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11842_ (.CLK(clk),
    .D(_00069_),
    .RESET_B(net247),
    .Q(\u_rf.reg0_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11843_ (.CLK(clk),
    .D(_00070_),
    .RESET_B(net250),
    .Q(\u_rf.reg0_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11844_ (.CLK(clk),
    .D(_00071_),
    .RESET_B(net234),
    .Q(\u_rf.reg0_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11845_ (.CLK(clk),
    .D(_00072_),
    .RESET_B(net314),
    .Q(\u_rf.reg0_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11846_ (.CLK(clk),
    .D(_00073_),
    .RESET_B(net317),
    .Q(\u_rf.reg0_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11847_ (.CLK(clk),
    .D(_00074_),
    .RESET_B(net247),
    .Q(\u_rf.reg0_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11848_ (.CLK(clk),
    .D(_00075_),
    .RESET_B(net202),
    .Q(\u_rf.reg0_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11849_ (.CLK(clk),
    .D(_00076_),
    .RESET_B(net211),
    .Q(\u_rf.reg0_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11850_ (.CLK(clk),
    .D(_00077_),
    .RESET_B(net288),
    .Q(\u_rf.reg0_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11851_ (.CLK(clk),
    .D(_00078_),
    .RESET_B(net280),
    .Q(\u_rf.reg0_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11852_ (.CLK(clk),
    .D(_00079_),
    .RESET_B(net257),
    .Q(\u_rf.reg0_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11853_ (.CLK(clk),
    .D(_00080_),
    .RESET_B(net208),
    .Q(\u_rf.reg0_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11854_ (.CLK(clk),
    .D(_00081_),
    .RESET_B(net244),
    .Q(\u_rf.reg0_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11855_ (.CLK(clk),
    .D(_00082_),
    .RESET_B(net215),
    .Q(\u_rf.reg0_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11856_ (.CLK(clk),
    .D(_00083_),
    .RESET_B(net256),
    .Q(\u_rf.reg0_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11857_ (.CLK(clk),
    .D(_00084_),
    .RESET_B(net276),
    .Q(\u_rf.reg0_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11858_ (.CLK(clk),
    .D(_00085_),
    .RESET_B(net276),
    .Q(\u_rf.reg0_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11859_ (.CLK(clk),
    .D(_00086_),
    .RESET_B(net284),
    .Q(\u_rf.reg0_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11860_ (.CLK(clk),
    .D(_00087_),
    .RESET_B(net277),
    .Q(\u_rf.reg0_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11861_ (.CLK(clk),
    .D(_00088_),
    .RESET_B(net355),
    .Q(\u_rf.reg0_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11862_ (.CLK(clk),
    .D(_00089_),
    .RESET_B(net269),
    .Q(\u_rf.reg0_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11863_ (.CLK(clk),
    .D(_00090_),
    .RESET_B(net296),
    .Q(\u_rf.reg0_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11864_ (.CLK(clk),
    .D(_00091_),
    .RESET_B(net307),
    .Q(\u_rf.reg0_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11865_ (.CLK(clk),
    .D(_00092_),
    .RESET_B(net358),
    .Q(\u_rf.reg0_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11866_ (.CLK(clk),
    .D(_00093_),
    .RESET_B(net355),
    .Q(\u_rf.reg0_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11867_ (.CLK(clk),
    .D(_00094_),
    .RESET_B(net343),
    .Q(\u_rf.reg0_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11868_ (.CLK(clk),
    .D(_00095_),
    .RESET_B(net340),
    .Q(\u_rf.reg0_q[31] ));
 sky130_fd_sc_hd__dfrtp_4 _11869_ (.CLK(clk),
    .D(\u_decod.dec0.operation_o[0] ),
    .RESET_B(net335),
    .Q(\u_decod.instr_operation_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11870_ (.CLK(clk),
    .D(\u_decod.dec0.operation_o[1] ),
    .RESET_B(net336),
    .Q(\u_decod.instr_operation_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11871_ (.CLK(clk),
    .D(\u_decod.dec0.operation_o[2] ),
    .RESET_B(net337),
    .Q(\u_decod.instr_operation_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11872_ (.CLK(clk),
    .D(\u_decod.dec0.operation_o[3] ),
    .RESET_B(net335),
    .Q(\u_decod.instr_operation_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11873_ (.CLK(clk),
    .D(\u_decod.dec0.operation_o[4] ),
    .RESET_B(net335),
    .Q(\u_decod.instr_operation_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11874_ (.CLK(clk),
    .D(\u_decod.dec0.jalr ),
    .RESET_B(net336),
    .Q(\u_decod.instr_operation_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11875_ (.CLK(clk),
    .D(\u_decod.dec0.unsign_extension ),
    .RESET_B(net332),
    .Q(\u_decod.unsign_ext_q_o ));
 sky130_fd_sc_hd__dfrtp_4 _11876_ (.CLK(clk),
    .D(\u_decod.dec0.access_size_o[0] ),
    .RESET_B(net335),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 _11877_ (.CLK(clk),
    .D(\u_decod.dec0.access_size_o[1] ),
    .RESET_B(net335),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _11878_ (.CLK(clk),
    .D(\u_decod.dec0.access_size_o[2] ),
    .RESET_B(net335),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _11879_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[0] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11880_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[1] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11881_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[2] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11882_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[3] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11883_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[4] ),
    .RESET_B(net335),
    .Q(\u_decod.rs2_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11884_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[5] ),
    .RESET_B(net322),
    .Q(\u_decod.rs2_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11885_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[6] ),
    .RESET_B(net322),
    .Q(\u_decod.rs2_data_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11886_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[7] ),
    .RESET_B(net322),
    .Q(\u_decod.rs2_data_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11887_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[8] ),
    .RESET_B(net322),
    .Q(\u_decod.rs2_data_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11888_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[9] ),
    .RESET_B(net334),
    .Q(\u_decod.rs2_data_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11889_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[10] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11890_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[11] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11891_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[12] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11892_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[13] ),
    .RESET_B(net329),
    .Q(\u_decod.rs2_data_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11893_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[14] ),
    .RESET_B(net332),
    .Q(\u_decod.rs2_data_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11894_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[15] ),
    .RESET_B(net333),
    .Q(\u_decod.rs2_data_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11895_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[16] ),
    .RESET_B(net332),
    .Q(\u_decod.rs2_data_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11896_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[17] ),
    .RESET_B(net332),
    .Q(\u_decod.rs2_data_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11897_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[18] ),
    .RESET_B(net333),
    .Q(\u_decod.rs2_data_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11898_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[19] ),
    .RESET_B(net333),
    .Q(\u_decod.rs2_data_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11899_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[20] ),
    .RESET_B(net345),
    .Q(\u_decod.rs2_data_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11900_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[21] ),
    .RESET_B(net345),
    .Q(\u_decod.rs2_data_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11901_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[22] ),
    .RESET_B(net345),
    .Q(\u_decod.rs2_data_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11902_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[23] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11903_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[24] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11904_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[25] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11905_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[26] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11906_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[27] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11907_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[28] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11908_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[29] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11909_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[30] ),
    .RESET_B(net347),
    .Q(\u_decod.rs2_data_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11910_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[31] ),
    .RESET_B(net345),
    .Q(\u_decod.rs2_data_q[31] ));
 sky130_fd_sc_hd__dfrtp_2 _11911_ (.CLK(clk),
    .D(\u_decod.rs2_data_nxt[32] ),
    .RESET_B(net345),
    .Q(\u_decod.rs2_data_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 _11912_ (.CLK(clk),
    .D(\u_decod.rs1_data[0] ),
    .RESET_B(net330),
    .Q(\u_decod.rs1_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11913_ (.CLK(clk),
    .D(\u_decod.rs1_data[1] ),
    .RESET_B(net336),
    .Q(\u_decod.rs1_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11914_ (.CLK(clk),
    .D(\u_decod.rs1_data[2] ),
    .RESET_B(net332),
    .Q(\u_decod.rs1_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11915_ (.CLK(clk),
    .D(\u_decod.rs1_data[3] ),
    .RESET_B(net336),
    .Q(\u_decod.rs1_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11916_ (.CLK(clk),
    .D(\u_decod.rs1_data[4] ),
    .RESET_B(net337),
    .Q(\u_decod.rs1_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11917_ (.CLK(clk),
    .D(\u_decod.rs1_data[5] ),
    .RESET_B(net332),
    .Q(\u_decod.rs1_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11918_ (.CLK(clk),
    .D(\u_decod.rs1_data[6] ),
    .RESET_B(net332),
    .Q(\u_decod.rs1_data_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11919_ (.CLK(clk),
    .D(\u_decod.rs1_data[7] ),
    .RESET_B(net337),
    .Q(\u_decod.rs1_data_q[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11920_ (.CLK(clk),
    .D(\u_decod.rs1_data[8] ),
    .RESET_B(net337),
    .Q(\u_decod.rs1_data_q[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11921_ (.CLK(clk),
    .D(\u_decod.rs1_data[9] ),
    .RESET_B(net337),
    .Q(\u_decod.rs1_data_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11922_ (.CLK(clk),
    .D(\u_decod.rs1_data[10] ),
    .RESET_B(net333),
    .Q(\u_decod.rs1_data_q[10] ));
 sky130_fd_sc_hd__dfrtp_4 _11923_ (.CLK(clk),
    .D(\u_decod.rs1_data[11] ),
    .RESET_B(net362),
    .Q(\u_decod.rs1_data_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11924_ (.CLK(clk),
    .D(\u_decod.rs1_data[12] ),
    .RESET_B(net362),
    .Q(\u_decod.rs1_data_q[12] ));
 sky130_fd_sc_hd__dfrtp_4 _11925_ (.CLK(clk),
    .D(\u_decod.rs1_data[13] ),
    .RESET_B(net360),
    .Q(\u_decod.rs1_data_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11926_ (.CLK(clk),
    .D(\u_decod.rs1_data[14] ),
    .RESET_B(net362),
    .Q(\u_decod.rs1_data_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11927_ (.CLK(clk),
    .D(\u_decod.rs1_data[15] ),
    .RESET_B(net362),
    .Q(\u_decod.rs1_data_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11928_ (.CLK(clk),
    .D(\u_decod.rs1_data[16] ),
    .RESET_B(net338),
    .Q(\u_decod.rs1_data_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11929_ (.CLK(clk),
    .D(\u_decod.rs1_data[17] ),
    .RESET_B(net338),
    .Q(\u_decod.rs1_data_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11930_ (.CLK(clk),
    .D(\u_decod.rs1_data[18] ),
    .RESET_B(net338),
    .Q(\u_decod.rs1_data_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11931_ (.CLK(clk),
    .D(\u_decod.rs1_data[19] ),
    .RESET_B(net338),
    .Q(\u_decod.rs1_data_q[19] ));
 sky130_fd_sc_hd__dfrtp_2 _11932_ (.CLK(clk),
    .D(\u_decod.rs1_data[20] ),
    .RESET_B(net371),
    .Q(\u_decod.rs1_data_q[20] ));
 sky130_fd_sc_hd__dfrtp_2 _11933_ (.CLK(clk),
    .D(\u_decod.rs1_data[21] ),
    .RESET_B(net371),
    .Q(\u_decod.rs1_data_q[21] ));
 sky130_fd_sc_hd__dfrtp_2 _11934_ (.CLK(clk),
    .D(\u_decod.rs1_data[22] ),
    .RESET_B(net370),
    .Q(\u_decod.rs1_data_q[22] ));
 sky130_fd_sc_hd__dfrtp_2 _11935_ (.CLK(clk),
    .D(\u_decod.rs1_data[23] ),
    .RESET_B(net370),
    .Q(\u_decod.rs1_data_q[23] ));
 sky130_fd_sc_hd__dfrtp_4 _11936_ (.CLK(clk),
    .D(\u_decod.rs1_data[24] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[24] ));
 sky130_fd_sc_hd__dfrtp_4 _11937_ (.CLK(clk),
    .D(\u_decod.rs1_data[25] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[25] ));
 sky130_fd_sc_hd__dfrtp_4 _11938_ (.CLK(clk),
    .D(\u_decod.rs1_data[26] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[26] ));
 sky130_fd_sc_hd__dfrtp_4 _11939_ (.CLK(clk),
    .D(\u_decod.rs1_data[27] ),
    .RESET_B(net358),
    .Q(\u_decod.rs1_data_q[27] ));
 sky130_fd_sc_hd__dfrtp_4 _11940_ (.CLK(clk),
    .D(\u_decod.rs1_data[28] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[28] ));
 sky130_fd_sc_hd__dfrtp_4 _11941_ (.CLK(clk),
    .D(\u_decod.rs1_data[29] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[29] ));
 sky130_fd_sc_hd__dfrtp_4 _11942_ (.CLK(clk),
    .D(\u_decod.rs1_data[30] ),
    .RESET_B(net357),
    .Q(\u_decod.rs1_data_q[30] ));
 sky130_fd_sc_hd__dfrtp_2 _11943_ (.CLK(clk),
    .D(\u_decod.rs1_data[31] ),
    .RESET_B(net362),
    .Q(\u_decod.rs1_data_q[31] ));
 sky130_fd_sc_hd__dfrtp_2 _11944_ (.CLK(clk),
    .D(\u_decod.rs1_data_nxt[32] ),
    .RESET_B(net345),
    .Q(\u_decod.rs1_data_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 _11945_ (.CLK(clk),
    .D(\u_decod.dec0.rd_v ),
    .RESET_B(net332),
    .Q(\u_decod.rd_v_q ));
 sky130_fd_sc_hd__dfrtp_4 _11946_ (.CLK(clk),
    .D(\u_decod.dec0.rd_o[0] ),
    .RESET_B(net328),
    .Q(\u_decod.exe_ff_rd_adr_q_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11947_ (.CLK(clk),
    .D(\u_decod.dec0.rd_o[1] ),
    .RESET_B(net331),
    .Q(\u_decod.exe_ff_rd_adr_q_i[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11948_ (.CLK(clk),
    .D(\u_decod.dec0.rd_o[2] ),
    .RESET_B(net325),
    .Q(\u_decod.exe_ff_rd_adr_q_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11949_ (.CLK(clk),
    .D(\u_decod.dec0.rd_o[3] ),
    .RESET_B(net331),
    .Q(\u_decod.exe_ff_rd_adr_q_i[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11950_ (.CLK(clk),
    .D(\u_decod.dec0.rd_o[4] ),
    .RESET_B(net325),
    .Q(\u_decod.exe_ff_rd_adr_q_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11951_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[0] ),
    .RESET_B(net332),
    .Q(\u_decod.pc_q_o[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11952_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[1] ),
    .RESET_B(net336),
    .Q(\u_decod.pc_q_o[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11953_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[2] ),
    .RESET_B(net338),
    .Q(\u_decod.pc_q_o[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11954_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[3] ),
    .RESET_B(net338),
    .Q(\u_decod.pc_q_o[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11955_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[4] ),
    .RESET_B(net338),
    .Q(\u_decod.pc_q_o[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11956_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[5] ),
    .RESET_B(net360),
    .Q(\u_decod.pc_q_o[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11957_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[6] ),
    .RESET_B(net338),
    .Q(\u_decod.pc_q_o[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11958_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[7] ),
    .RESET_B(net338),
    .Q(\u_decod.pc_q_o[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11959_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[8] ),
    .RESET_B(net374),
    .Q(\u_decod.pc_q_o[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11960_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[9] ),
    .RESET_B(net362),
    .Q(\u_decod.pc_q_o[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11961_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[10] ),
    .RESET_B(net360),
    .Q(\u_decod.pc_q_o[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11962_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[11] ),
    .RESET_B(net362),
    .Q(\u_decod.pc_q_o[11] ));
 sky130_fd_sc_hd__dfrtp_4 _11963_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[12] ),
    .RESET_B(net366),
    .Q(\u_decod.pc_q_o[12] ));
 sky130_fd_sc_hd__dfrtp_4 _11964_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[13] ),
    .RESET_B(net366),
    .Q(\u_decod.pc_q_o[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11965_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[14] ),
    .RESET_B(net366),
    .Q(\u_decod.pc_q_o[14] ));
 sky130_fd_sc_hd__dfrtp_2 _11966_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[15] ),
    .RESET_B(net361),
    .Q(\u_decod.pc_q_o[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11967_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[16] ),
    .RESET_B(net365),
    .Q(\u_decod.pc_q_o[16] ));
 sky130_fd_sc_hd__dfrtp_2 _11968_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[17] ),
    .RESET_B(net365),
    .Q(\u_decod.pc_q_o[17] ));
 sky130_fd_sc_hd__dfrtp_2 _11969_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[18] ),
    .RESET_B(net372),
    .Q(\u_decod.pc_q_o[18] ));
 sky130_fd_sc_hd__dfrtp_2 _11970_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[19] ),
    .RESET_B(net372),
    .Q(\u_decod.pc_q_o[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11971_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[20] ),
    .RESET_B(net370),
    .Q(\u_decod.pc_q_o[20] ));
 sky130_fd_sc_hd__dfrtp_4 _11972_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[21] ),
    .RESET_B(net370),
    .Q(\u_decod.pc_q_o[21] ));
 sky130_fd_sc_hd__dfrtp_4 _11973_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[22] ),
    .RESET_B(net370),
    .Q(\u_decod.pc_q_o[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11974_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[23] ),
    .RESET_B(net371),
    .Q(\u_decod.pc_q_o[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11975_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[24] ),
    .RESET_B(net368),
    .Q(\u_decod.pc_q_o[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11976_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[25] ),
    .RESET_B(net368),
    .Q(\u_decod.pc_q_o[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11977_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[26] ),
    .RESET_B(net369),
    .Q(\u_decod.pc_q_o[26] ));
 sky130_fd_sc_hd__dfrtp_2 _11978_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[27] ),
    .RESET_B(net369),
    .Q(\u_decod.pc_q_o[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11979_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[28] ),
    .RESET_B(net368),
    .Q(\u_decod.pc_q_o[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11980_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[29] ),
    .RESET_B(net357),
    .Q(\u_decod.pc_q_o[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11981_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[30] ),
    .RESET_B(net357),
    .Q(\u_decod.pc_q_o[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11982_ (.CLK(clk),
    .D(\u_decod.pc0_q_i[31] ),
    .RESET_B(net347),
    .Q(\u_decod.pc_q_o[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11983_ (.CLK(clk),
    .D(\u_decod.dec0.is_arithm ),
    .RESET_B(net335),
    .Q(\u_decod.instr_unit_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11984_ (.CLK(clk),
    .D(\u_decod.dec0.is_shift ),
    .RESET_B(net335),
    .Q(\u_decod.instr_unit_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11985_ (.CLK(clk),
    .D(\u_decod.dec0.is_branch ),
    .RESET_B(net336),
    .Q(\u_decod.instr_unit_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11986_ (.CLK(clk),
    .D(\u_decod.dec0.unit_o[3] ),
    .RESET_B(net335),
    .Q(\u_decod.instr_unit_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11987_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[0] ),
    .RESET_B(net360),
    .Q(\u_exe.pc_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11988_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[1] ),
    .RESET_B(net360),
    .Q(\u_exe.pc_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11989_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[2] ),
    .RESET_B(net361),
    .Q(\u_exe.pc_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11990_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[3] ),
    .RESET_B(net361),
    .Q(\u_exe.pc_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11991_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[4] ),
    .RESET_B(net361),
    .Q(\u_exe.pc_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11992_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[5] ),
    .RESET_B(net362),
    .Q(\u_exe.pc_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11993_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[6] ),
    .RESET_B(net364),
    .Q(\u_exe.pc_data_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11994_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[7] ),
    .RESET_B(net363),
    .Q(\u_exe.pc_data_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11995_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[8] ),
    .RESET_B(net363),
    .Q(\u_exe.pc_data_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11996_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[9] ),
    .RESET_B(net363),
    .Q(\u_exe.pc_data_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11997_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[10] ),
    .RESET_B(net364),
    .Q(\u_exe.pc_data_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11998_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[11] ),
    .RESET_B(net364),
    .Q(\u_exe.pc_data_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11999_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[12] ),
    .RESET_B(net364),
    .Q(\u_exe.pc_data_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12000_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[13] ),
    .RESET_B(net365),
    .Q(\u_exe.pc_data_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12001_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[14] ),
    .RESET_B(net366),
    .Q(\u_exe.pc_data_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12002_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[15] ),
    .RESET_B(net366),
    .Q(\u_exe.pc_data_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12003_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[16] ),
    .RESET_B(net366),
    .Q(\u_exe.pc_data_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12004_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[17] ),
    .RESET_B(net365),
    .Q(\u_exe.pc_data_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12005_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[18] ),
    .RESET_B(net370),
    .Q(\u_exe.pc_data_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12006_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[19] ),
    .RESET_B(net372),
    .Q(\u_exe.pc_data_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12007_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[20] ),
    .RESET_B(net372),
    .Q(\u_exe.pc_data_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12008_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[21] ),
    .RESET_B(net371),
    .Q(\u_exe.pc_data_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12009_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[22] ),
    .RESET_B(net371),
    .Q(\u_exe.pc_data_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12010_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[23] ),
    .RESET_B(net371),
    .Q(\u_exe.pc_data_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12011_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[24] ),
    .RESET_B(net369),
    .Q(\u_exe.pc_data_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12012_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[25] ),
    .RESET_B(net368),
    .Q(\u_exe.pc_data_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12013_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[26] ),
    .RESET_B(net369),
    .Q(\u_exe.pc_data_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12014_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[27] ),
    .RESET_B(net369),
    .Q(\u_exe.pc_data_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12015_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[28] ),
    .RESET_B(net368),
    .Q(\u_exe.pc_data_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12016_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[29] ),
    .RESET_B(net368),
    .Q(\u_exe.pc_data_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12017_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[30] ),
    .RESET_B(net368),
    .Q(\u_exe.pc_data_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12018_ (.CLK(clk),
    .D(\u_exe.bu_pc_res[31] ),
    .RESET_B(net367),
    .Q(\u_exe.pc_data_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12019_ (.CLK(clk),
    .D(\u_decod.flush_v ),
    .RESET_B(net332),
    .Q(\u_exe.flush_v_dly1_q ));
 sky130_fd_sc_hd__dfrtp_4 _12020_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[0] ),
    .RESET_B(net330),
    .Q(\u_decod.rf_ff_res_data_i[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12021_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[1] ),
    .RESET_B(net328),
    .Q(\u_decod.rf_ff_res_data_i[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12022_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[2] ),
    .RESET_B(net331),
    .Q(\u_decod.rf_ff_res_data_i[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12023_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[3] ),
    .RESET_B(net328),
    .Q(\u_decod.rf_ff_res_data_i[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12024_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[4] ),
    .RESET_B(net322),
    .Q(\u_decod.rf_ff_res_data_i[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12025_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[5] ),
    .RESET_B(net330),
    .Q(\u_decod.rf_ff_res_data_i[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12026_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[6] ),
    .RESET_B(net331),
    .Q(\u_decod.rf_ff_res_data_i[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12027_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[7] ),
    .RESET_B(net322),
    .Q(\u_decod.rf_ff_res_data_i[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12028_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[8] ),
    .RESET_B(net321),
    .Q(\u_decod.rf_ff_res_data_i[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12029_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[9] ),
    .RESET_B(net322),
    .Q(\u_decod.rf_ff_res_data_i[9] ));
 sky130_fd_sc_hd__dfrtp_4 _12030_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[10] ),
    .RESET_B(net328),
    .Q(\u_decod.rf_ff_res_data_i[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12031_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[11] ),
    .RESET_B(net328),
    .Q(\u_decod.rf_ff_res_data_i[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12032_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[12] ),
    .RESET_B(net330),
    .Q(\u_decod.rf_ff_res_data_i[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12033_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[13] ),
    .RESET_B(net344),
    .Q(\u_decod.rf_ff_res_data_i[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12034_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[14] ),
    .RESET_B(net344),
    .Q(\u_decod.rf_ff_res_data_i[14] ));
 sky130_fd_sc_hd__dfrtp_4 _12035_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[15] ),
    .RESET_B(net344),
    .Q(\u_decod.rf_ff_res_data_i[15] ));
 sky130_fd_sc_hd__dfrtp_4 _12036_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[16] ),
    .RESET_B(net331),
    .Q(\u_decod.rf_ff_res_data_i[16] ));
 sky130_fd_sc_hd__dfrtp_4 _12037_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[17] ),
    .RESET_B(net331),
    .Q(\u_decod.rf_ff_res_data_i[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12038_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[18] ),
    .RESET_B(net331),
    .Q(\u_decod.rf_ff_res_data_i[18] ));
 sky130_fd_sc_hd__dfrtp_4 _12039_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[19] ),
    .RESET_B(net333),
    .Q(\u_decod.rf_ff_res_data_i[19] ));
 sky130_fd_sc_hd__dfrtp_4 _12040_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[20] ),
    .RESET_B(net355),
    .Q(\u_decod.rf_ff_res_data_i[20] ));
 sky130_fd_sc_hd__dfrtp_4 _12041_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[21] ),
    .RESET_B(net355),
    .Q(\u_decod.rf_ff_res_data_i[21] ));
 sky130_fd_sc_hd__dfrtp_4 _12042_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[22] ),
    .RESET_B(net346),
    .Q(\u_decod.rf_ff_res_data_i[22] ));
 sky130_fd_sc_hd__dfrtp_4 _12043_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[23] ),
    .RESET_B(net358),
    .Q(\u_decod.rf_ff_res_data_i[23] ));
 sky130_fd_sc_hd__dfrtp_2 _12044_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[24] ),
    .RESET_B(net356),
    .Q(\u_decod.rf_ff_res_data_i[24] ));
 sky130_fd_sc_hd__dfrtp_4 _12045_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[25] ),
    .RESET_B(net346),
    .Q(\u_decod.rf_ff_res_data_i[25] ));
 sky130_fd_sc_hd__dfrtp_4 _12046_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[26] ),
    .RESET_B(net356),
    .Q(\u_decod.rf_ff_res_data_i[26] ));
 sky130_fd_sc_hd__dfrtp_4 _12047_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[27] ),
    .RESET_B(net358),
    .Q(\u_decod.rf_ff_res_data_i[27] ));
 sky130_fd_sc_hd__dfrtp_4 _12048_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[28] ),
    .RESET_B(net355),
    .Q(\u_decod.rf_ff_res_data_i[28] ));
 sky130_fd_sc_hd__dfrtp_2 _12049_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[29] ),
    .RESET_B(net357),
    .Q(\u_decod.rf_ff_res_data_i[29] ));
 sky130_fd_sc_hd__dfrtp_2 _12050_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[30] ),
    .RESET_B(net346),
    .Q(\u_decod.rf_ff_res_data_i[30] ));
 sky130_fd_sc_hd__dfrtp_2 _12051_ (.CLK(clk),
    .D(\u_decod.exe_ff_res_data_i[31] ),
    .RESET_B(net344),
    .Q(\u_decod.rf_ff_res_data_i[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12052_ (.CLK(clk),
    .D(\u_decod.exe_ff_write_v_q_i ),
    .RESET_B(net333),
    .Q(\u_decod.rf_write_v_q_i ));
 sky130_fd_sc_hd__dfrtp_4 _12053_ (.CLK(clk),
    .D(\u_decod.exe_ff_rd_adr_q_i[0] ),
    .RESET_B(net325),
    .Q(\u_decod.rf_ff_rd_adr_q_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12054_ (.CLK(clk),
    .D(\u_decod.exe_ff_rd_adr_q_i[1] ),
    .RESET_B(net333),
    .Q(\u_decod.rf_ff_rd_adr_q_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12055_ (.CLK(clk),
    .D(\u_decod.exe_ff_rd_adr_q_i[2] ),
    .RESET_B(net325),
    .Q(\u_decod.rf_ff_rd_adr_q_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12056_ (.CLK(clk),
    .D(\u_decod.exe_ff_rd_adr_q_i[3] ),
    .RESET_B(net333),
    .Q(\u_decod.rf_ff_rd_adr_q_i[3] ));
 sky130_fd_sc_hd__dfrtp_2 _12057_ (.CLK(clk),
    .D(\u_decod.exe_ff_rd_adr_q_i[4] ),
    .RESET_B(net327),
    .Q(\u_decod.rf_ff_rd_adr_q_i[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12058_ (.CLK(clk),
    .D(\u_exe.branch_v ),
    .RESET_B(net361),
    .Q(\u_decod.flush_v ));
 sky130_fd_sc_hd__dfrtp_1 _12059_ (.CLK(clk),
    .D(_00096_),
    .RESET_B(net221),
    .Q(\u_rf.reg3_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12060_ (.CLK(clk),
    .D(_00097_),
    .RESET_B(net236),
    .Q(\u_rf.reg3_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12061_ (.CLK(clk),
    .D(_00098_),
    .RESET_B(net250),
    .Q(\u_rf.reg3_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12062_ (.CLK(clk),
    .D(_00099_),
    .RESET_B(net209),
    .Q(\u_rf.reg3_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12063_ (.CLK(clk),
    .D(_00100_),
    .RESET_B(net227),
    .Q(\u_rf.reg3_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12064_ (.CLK(clk),
    .D(_00101_),
    .RESET_B(net247),
    .Q(\u_rf.reg3_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12065_ (.CLK(clk),
    .D(_00102_),
    .RESET_B(net251),
    .Q(\u_rf.reg3_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12066_ (.CLK(clk),
    .D(_00103_),
    .RESET_B(net229),
    .Q(\u_rf.reg3_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12067_ (.CLK(clk),
    .D(_00104_),
    .RESET_B(net312),
    .Q(\u_rf.reg3_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12068_ (.CLK(clk),
    .D(_00105_),
    .RESET_B(net312),
    .Q(\u_rf.reg3_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12069_ (.CLK(clk),
    .D(_00106_),
    .RESET_B(net239),
    .Q(\u_rf.reg3_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12070_ (.CLK(clk),
    .D(_00107_),
    .RESET_B(net202),
    .Q(\u_rf.reg3_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12071_ (.CLK(clk),
    .D(_00108_),
    .RESET_B(net211),
    .Q(\u_rf.reg3_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12072_ (.CLK(clk),
    .D(_00109_),
    .RESET_B(net288),
    .Q(\u_rf.reg3_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12073_ (.CLK(clk),
    .D(_00110_),
    .RESET_B(net265),
    .Q(\u_rf.reg3_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12074_ (.CLK(clk),
    .D(_00111_),
    .RESET_B(net257),
    .Q(\u_rf.reg3_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12075_ (.CLK(clk),
    .D(_00112_),
    .RESET_B(net208),
    .Q(\u_rf.reg3_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12076_ (.CLK(clk),
    .D(_00113_),
    .RESET_B(net266),
    .Q(\u_rf.reg3_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12077_ (.CLK(clk),
    .D(_00114_),
    .RESET_B(net215),
    .Q(\u_rf.reg3_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12078_ (.CLK(clk),
    .D(_00115_),
    .RESET_B(net256),
    .Q(\u_rf.reg3_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12079_ (.CLK(clk),
    .D(_00116_),
    .RESET_B(net272),
    .Q(\u_rf.reg3_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12080_ (.CLK(clk),
    .D(_00117_),
    .RESET_B(net271),
    .Q(\u_rf.reg3_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12081_ (.CLK(clk),
    .D(_00118_),
    .RESET_B(net294),
    .Q(\u_rf.reg3_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12082_ (.CLK(clk),
    .D(_00119_),
    .RESET_B(net277),
    .Q(\u_rf.reg3_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12083_ (.CLK(clk),
    .D(_00120_),
    .RESET_B(net304),
    .Q(\u_rf.reg3_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12084_ (.CLK(clk),
    .D(_00121_),
    .RESET_B(net269),
    .Q(\u_rf.reg3_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12085_ (.CLK(clk),
    .D(_00122_),
    .RESET_B(net300),
    .Q(\u_rf.reg3_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12086_ (.CLK(clk),
    .D(_00123_),
    .RESET_B(net306),
    .Q(\u_rf.reg3_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12087_ (.CLK(clk),
    .D(_00124_),
    .RESET_B(net308),
    .Q(\u_rf.reg3_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12088_ (.CLK(clk),
    .D(_00125_),
    .RESET_B(net292),
    .Q(\u_rf.reg3_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12089_ (.CLK(clk),
    .D(_00126_),
    .RESET_B(net291),
    .Q(\u_rf.reg3_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12090_ (.CLK(clk),
    .D(_00127_),
    .RESET_B(net289),
    .Q(\u_rf.reg3_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12091_ (.CLK(clk),
    .D(_00128_),
    .RESET_B(net222),
    .Q(\u_rf.reg4_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12092_ (.CLK(clk),
    .D(_00129_),
    .RESET_B(net234),
    .Q(\u_rf.reg4_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12093_ (.CLK(clk),
    .D(_00130_),
    .RESET_B(net245),
    .Q(\u_rf.reg4_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12094_ (.CLK(clk),
    .D(_00131_),
    .RESET_B(net209),
    .Q(\u_rf.reg4_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12095_ (.CLK(clk),
    .D(_00132_),
    .RESET_B(net206),
    .Q(\u_rf.reg4_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12096_ (.CLK(clk),
    .D(_00133_),
    .RESET_B(net323),
    .Q(\u_rf.reg4_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12097_ (.CLK(clk),
    .D(_00134_),
    .RESET_B(net250),
    .Q(\u_rf.reg4_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12098_ (.CLK(clk),
    .D(_00135_),
    .RESET_B(net229),
    .Q(\u_rf.reg4_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12099_ (.CLK(clk),
    .D(_00136_),
    .RESET_B(net314),
    .Q(\u_rf.reg4_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12100_ (.CLK(clk),
    .D(_00137_),
    .RESET_B(net314),
    .Q(\u_rf.reg4_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12101_ (.CLK(clk),
    .D(_00138_),
    .RESET_B(net239),
    .Q(\u_rf.reg4_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12102_ (.CLK(clk),
    .D(_00139_),
    .RESET_B(net202),
    .Q(\u_rf.reg4_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12103_ (.CLK(clk),
    .D(_00140_),
    .RESET_B(net212),
    .Q(\u_rf.reg4_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12104_ (.CLK(clk),
    .D(_00141_),
    .RESET_B(net281),
    .Q(\u_rf.reg4_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12105_ (.CLK(clk),
    .D(_00142_),
    .RESET_B(net284),
    .Q(\u_rf.reg4_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12106_ (.CLK(clk),
    .D(_00143_),
    .RESET_B(net261),
    .Q(\u_rf.reg4_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12107_ (.CLK(clk),
    .D(_00144_),
    .RESET_B(net208),
    .Q(\u_rf.reg4_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12108_ (.CLK(clk),
    .D(_00145_),
    .RESET_B(net226),
    .Q(\u_rf.reg4_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12109_ (.CLK(clk),
    .D(_00146_),
    .RESET_B(net215),
    .Q(\u_rf.reg4_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12110_ (.CLK(clk),
    .D(_00147_),
    .RESET_B(net256),
    .Q(\u_rf.reg4_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12111_ (.CLK(clk),
    .D(_00148_),
    .RESET_B(net275),
    .Q(\u_rf.reg4_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12112_ (.CLK(clk),
    .D(_00149_),
    .RESET_B(net284),
    .Q(\u_rf.reg4_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12113_ (.CLK(clk),
    .D(_00150_),
    .RESET_B(net296),
    .Q(\u_rf.reg4_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12114_ (.CLK(clk),
    .D(_00151_),
    .RESET_B(net298),
    .Q(\u_rf.reg4_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12115_ (.CLK(clk),
    .D(_00152_),
    .RESET_B(net304),
    .Q(\u_rf.reg4_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12116_ (.CLK(clk),
    .D(_00153_),
    .RESET_B(net267),
    .Q(\u_rf.reg4_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12117_ (.CLK(clk),
    .D(_00154_),
    .RESET_B(net294),
    .Q(\u_rf.reg4_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12118_ (.CLK(clk),
    .D(_00155_),
    .RESET_B(net308),
    .Q(\u_rf.reg4_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12119_ (.CLK(clk),
    .D(_00156_),
    .RESET_B(net358),
    .Q(\u_rf.reg4_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12120_ (.CLK(clk),
    .D(_00157_),
    .RESET_B(net346),
    .Q(\u_rf.reg4_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12121_ (.CLK(clk),
    .D(_00158_),
    .RESET_B(net291),
    .Q(\u_rf.reg4_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12122_ (.CLK(clk),
    .D(_00159_),
    .RESET_B(net289),
    .Q(\u_rf.reg4_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12123_ (.CLK(clk),
    .D(_00160_),
    .RESET_B(net224),
    .Q(\u_rf.reg5_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12124_ (.CLK(clk),
    .D(_00161_),
    .RESET_B(net236),
    .Q(\u_rf.reg5_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12125_ (.CLK(clk),
    .D(_00162_),
    .RESET_B(net244),
    .Q(\u_rf.reg5_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12126_ (.CLK(clk),
    .D(_00163_),
    .RESET_B(net232),
    .Q(\u_rf.reg5_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12127_ (.CLK(clk),
    .D(_00164_),
    .RESET_B(net206),
    .Q(\u_rf.reg5_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12128_ (.CLK(clk),
    .D(_00165_),
    .RESET_B(net247),
    .Q(\u_rf.reg5_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12129_ (.CLK(clk),
    .D(_00166_),
    .RESET_B(net326),
    .Q(\u_rf.reg5_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12130_ (.CLK(clk),
    .D(_00167_),
    .RESET_B(net229),
    .Q(\u_rf.reg5_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12131_ (.CLK(clk),
    .D(_00168_),
    .RESET_B(net312),
    .Q(\u_rf.reg5_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12132_ (.CLK(clk),
    .D(_00169_),
    .RESET_B(net316),
    .Q(\u_rf.reg5_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12133_ (.CLK(clk),
    .D(_00170_),
    .RESET_B(net231),
    .Q(\u_rf.reg5_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12134_ (.CLK(clk),
    .D(_00171_),
    .RESET_B(net202),
    .Q(\u_rf.reg5_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12135_ (.CLK(clk),
    .D(_00172_),
    .RESET_B(net211),
    .Q(\u_rf.reg5_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12136_ (.CLK(clk),
    .D(_00173_),
    .RESET_B(net288),
    .Q(\u_rf.reg5_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12137_ (.CLK(clk),
    .D(_00174_),
    .RESET_B(net265),
    .Q(\u_rf.reg5_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12138_ (.CLK(clk),
    .D(_00175_),
    .RESET_B(net257),
    .Q(\u_rf.reg5_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12139_ (.CLK(clk),
    .D(_00176_),
    .RESET_B(net208),
    .Q(\u_rf.reg5_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12140_ (.CLK(clk),
    .D(_00177_),
    .RESET_B(net266),
    .Q(\u_rf.reg5_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12141_ (.CLK(clk),
    .D(_00178_),
    .RESET_B(net215),
    .Q(\u_rf.reg5_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12142_ (.CLK(clk),
    .D(_00179_),
    .RESET_B(net216),
    .Q(\u_rf.reg5_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12143_ (.CLK(clk),
    .D(_00180_),
    .RESET_B(net274),
    .Q(\u_rf.reg5_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12144_ (.CLK(clk),
    .D(_00181_),
    .RESET_B(net263),
    .Q(\u_rf.reg5_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12145_ (.CLK(clk),
    .D(_00182_),
    .RESET_B(net284),
    .Q(\u_rf.reg5_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12146_ (.CLK(clk),
    .D(_00183_),
    .RESET_B(net277),
    .Q(\u_rf.reg5_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12147_ (.CLK(clk),
    .D(_00184_),
    .RESET_B(net356),
    .Q(\u_rf.reg5_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12148_ (.CLK(clk),
    .D(_00185_),
    .RESET_B(net262),
    .Q(\u_rf.reg5_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12149_ (.CLK(clk),
    .D(_00186_),
    .RESET_B(net298),
    .Q(\u_rf.reg5_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12150_ (.CLK(clk),
    .D(_00187_),
    .RESET_B(net300),
    .Q(\u_rf.reg5_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12151_ (.CLK(clk),
    .D(_00188_),
    .RESET_B(net354),
    .Q(\u_rf.reg5_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12152_ (.CLK(clk),
    .D(_00189_),
    .RESET_B(net349),
    .Q(\u_rf.reg5_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12153_ (.CLK(clk),
    .D(_00190_),
    .RESET_B(net291),
    .Q(\u_rf.reg5_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12154_ (.CLK(clk),
    .D(_00191_),
    .RESET_B(net292),
    .Q(\u_rf.reg5_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12155_ (.CLK(clk),
    .D(_00192_),
    .RESET_B(net224),
    .Q(\u_rf.reg6_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12156_ (.CLK(clk),
    .D(_00193_),
    .RESET_B(net239),
    .Q(\u_rf.reg6_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12157_ (.CLK(clk),
    .D(_00194_),
    .RESET_B(net244),
    .Q(\u_rf.reg6_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12158_ (.CLK(clk),
    .D(_00195_),
    .RESET_B(net209),
    .Q(\u_rf.reg6_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12159_ (.CLK(clk),
    .D(_00196_),
    .RESET_B(net206),
    .Q(\u_rf.reg6_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12160_ (.CLK(clk),
    .D(_00197_),
    .RESET_B(net323),
    .Q(\u_rf.reg6_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12161_ (.CLK(clk),
    .D(_00198_),
    .RESET_B(net326),
    .Q(\u_rf.reg6_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12162_ (.CLK(clk),
    .D(_00199_),
    .RESET_B(net229),
    .Q(\u_rf.reg6_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12163_ (.CLK(clk),
    .D(_00200_),
    .RESET_B(net319),
    .Q(\u_rf.reg6_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12164_ (.CLK(clk),
    .D(_00201_),
    .RESET_B(net319),
    .Q(\u_rf.reg6_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12165_ (.CLK(clk),
    .D(_00202_),
    .RESET_B(net241),
    .Q(\u_rf.reg6_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12166_ (.CLK(clk),
    .D(_00203_),
    .RESET_B(net202),
    .Q(\u_rf.reg6_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12167_ (.CLK(clk),
    .D(_00204_),
    .RESET_B(net211),
    .Q(\u_rf.reg6_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12168_ (.CLK(clk),
    .D(_00205_),
    .RESET_B(net288),
    .Q(\u_rf.reg6_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12169_ (.CLK(clk),
    .D(_00206_),
    .RESET_B(net267),
    .Q(\u_rf.reg6_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12170_ (.CLK(clk),
    .D(_00207_),
    .RESET_B(net261),
    .Q(\u_rf.reg6_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12171_ (.CLK(clk),
    .D(_00208_),
    .RESET_B(net208),
    .Q(\u_rf.reg6_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12172_ (.CLK(clk),
    .D(_00209_),
    .RESET_B(net266),
    .Q(\u_rf.reg6_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12173_ (.CLK(clk),
    .D(_00210_),
    .RESET_B(net216),
    .Q(\u_rf.reg6_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12174_ (.CLK(clk),
    .D(_00211_),
    .RESET_B(net256),
    .Q(\u_rf.reg6_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12175_ (.CLK(clk),
    .D(_00212_),
    .RESET_B(net272),
    .Q(\u_rf.reg6_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12176_ (.CLK(clk),
    .D(_00213_),
    .RESET_B(net271),
    .Q(\u_rf.reg6_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12177_ (.CLK(clk),
    .D(_00214_),
    .RESET_B(net293),
    .Q(\u_rf.reg6_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12178_ (.CLK(clk),
    .D(_00215_),
    .RESET_B(net278),
    .Q(\u_rf.reg6_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12179_ (.CLK(clk),
    .D(_00216_),
    .RESET_B(net302),
    .Q(\u_rf.reg6_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12180_ (.CLK(clk),
    .D(_00217_),
    .RESET_B(net262),
    .Q(\u_rf.reg6_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12181_ (.CLK(clk),
    .D(_00218_),
    .RESET_B(net298),
    .Q(\u_rf.reg6_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12182_ (.CLK(clk),
    .D(_00219_),
    .RESET_B(net306),
    .Q(\u_rf.reg6_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12183_ (.CLK(clk),
    .D(_00220_),
    .RESET_B(net352),
    .Q(\u_rf.reg6_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12184_ (.CLK(clk),
    .D(_00221_),
    .RESET_B(net304),
    .Q(\u_rf.reg6_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12185_ (.CLK(clk),
    .D(_00222_),
    .RESET_B(net291),
    .Q(\u_rf.reg6_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12186_ (.CLK(clk),
    .D(_00223_),
    .RESET_B(net341),
    .Q(\u_rf.reg6_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12187_ (.CLK(clk),
    .D(_00224_),
    .RESET_B(net244),
    .Q(\u_rf.reg7_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12188_ (.CLK(clk),
    .D(_00225_),
    .RESET_B(net237),
    .Q(\u_rf.reg7_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12189_ (.CLK(clk),
    .D(_00226_),
    .RESET_B(net245),
    .Q(\u_rf.reg7_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12190_ (.CLK(clk),
    .D(_00227_),
    .RESET_B(net232),
    .Q(\u_rf.reg7_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12191_ (.CLK(clk),
    .D(_00228_),
    .RESET_B(net228),
    .Q(\u_rf.reg7_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12192_ (.CLK(clk),
    .D(_00229_),
    .RESET_B(net324),
    .Q(\u_rf.reg7_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12193_ (.CLK(clk),
    .D(_00230_),
    .RESET_B(net325),
    .Q(\u_rf.reg7_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12194_ (.CLK(clk),
    .D(_00231_),
    .RESET_B(net235),
    .Q(\u_rf.reg7_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12195_ (.CLK(clk),
    .D(_00232_),
    .RESET_B(net313),
    .Q(\u_rf.reg7_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12196_ (.CLK(clk),
    .D(_00233_),
    .RESET_B(net313),
    .Q(\u_rf.reg7_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12197_ (.CLK(clk),
    .D(_00234_),
    .RESET_B(net248),
    .Q(\u_rf.reg7_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12198_ (.CLK(clk),
    .D(_00235_),
    .RESET_B(net203),
    .Q(\u_rf.reg7_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12199_ (.CLK(clk),
    .D(_00236_),
    .RESET_B(net213),
    .Q(\u_rf.reg7_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12200_ (.CLK(clk),
    .D(_00237_),
    .RESET_B(net289),
    .Q(\u_rf.reg7_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12201_ (.CLK(clk),
    .D(_00238_),
    .RESET_B(net281),
    .Q(\u_rf.reg7_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12202_ (.CLK(clk),
    .D(_00239_),
    .RESET_B(net266),
    .Q(\u_rf.reg7_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12203_ (.CLK(clk),
    .D(_00240_),
    .RESET_B(net221),
    .Q(\u_rf.reg7_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12204_ (.CLK(clk),
    .D(_00241_),
    .RESET_B(net281),
    .Q(\u_rf.reg7_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12205_ (.CLK(clk),
    .D(_00242_),
    .RESET_B(net217),
    .Q(\u_rf.reg7_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12206_ (.CLK(clk),
    .D(_00243_),
    .RESET_B(net258),
    .Q(\u_rf.reg7_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12207_ (.CLK(clk),
    .D(_00244_),
    .RESET_B(net273),
    .Q(\u_rf.reg7_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12208_ (.CLK(clk),
    .D(_00245_),
    .RESET_B(net273),
    .Q(\u_rf.reg7_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12209_ (.CLK(clk),
    .D(_00246_),
    .RESET_B(net302),
    .Q(\u_rf.reg7_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12210_ (.CLK(clk),
    .D(_00247_),
    .RESET_B(net277),
    .Q(\u_rf.reg7_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12211_ (.CLK(clk),
    .D(_00248_),
    .RESET_B(net349),
    .Q(\u_rf.reg7_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12212_ (.CLK(clk),
    .D(_00249_),
    .RESET_B(net261),
    .Q(\u_rf.reg7_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12213_ (.CLK(clk),
    .D(_00250_),
    .RESET_B(net300),
    .Q(\u_rf.reg7_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12214_ (.CLK(clk),
    .D(_00251_),
    .RESET_B(net306),
    .Q(\u_rf.reg7_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12215_ (.CLK(clk),
    .D(_00252_),
    .RESET_B(net353),
    .Q(\u_rf.reg7_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12216_ (.CLK(clk),
    .D(_00253_),
    .RESET_B(net292),
    .Q(\u_rf.reg7_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12217_ (.CLK(clk),
    .D(_00254_),
    .RESET_B(net292),
    .Q(\u_rf.reg7_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12218_ (.CLK(clk),
    .D(_00255_),
    .RESET_B(net339),
    .Q(\u_rf.reg7_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12219_ (.CLK(clk),
    .D(_00256_),
    .RESET_B(net243),
    .Q(\u_rf.reg8_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12220_ (.CLK(clk),
    .D(_00257_),
    .RESET_B(net236),
    .Q(\u_rf.reg8_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12221_ (.CLK(clk),
    .D(_00258_),
    .RESET_B(net250),
    .Q(\u_rf.reg8_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12222_ (.CLK(clk),
    .D(_00259_),
    .RESET_B(net243),
    .Q(\u_rf.reg8_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12223_ (.CLK(clk),
    .D(_00260_),
    .RESET_B(net227),
    .Q(\u_rf.reg8_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12224_ (.CLK(clk),
    .D(_00261_),
    .RESET_B(net248),
    .Q(\u_rf.reg8_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12225_ (.CLK(clk),
    .D(_00262_),
    .RESET_B(net251),
    .Q(\u_rf.reg8_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12226_ (.CLK(clk),
    .D(_00263_),
    .RESET_B(net229),
    .Q(\u_rf.reg8_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12227_ (.CLK(clk),
    .D(_00264_),
    .RESET_B(net314),
    .Q(\u_rf.reg8_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12228_ (.CLK(clk),
    .D(_00265_),
    .RESET_B(net314),
    .Q(\u_rf.reg8_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12229_ (.CLK(clk),
    .D(_00266_),
    .RESET_B(net239),
    .Q(\u_rf.reg8_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12230_ (.CLK(clk),
    .D(_00267_),
    .RESET_B(net202),
    .Q(\u_rf.reg8_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12231_ (.CLK(clk),
    .D(_00268_),
    .RESET_B(net211),
    .Q(\u_rf.reg8_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12232_ (.CLK(clk),
    .D(_00269_),
    .RESET_B(net281),
    .Q(\u_rf.reg8_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12233_ (.CLK(clk),
    .D(_00270_),
    .RESET_B(net266),
    .Q(\u_rf.reg8_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12234_ (.CLK(clk),
    .D(_00271_),
    .RESET_B(net257),
    .Q(\u_rf.reg8_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12235_ (.CLK(clk),
    .D(_00272_),
    .RESET_B(net221),
    .Q(\u_rf.reg8_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12236_ (.CLK(clk),
    .D(_00273_),
    .RESET_B(net265),
    .Q(\u_rf.reg8_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12237_ (.CLK(clk),
    .D(_00274_),
    .RESET_B(net215),
    .Q(\u_rf.reg8_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12238_ (.CLK(clk),
    .D(_00275_),
    .RESET_B(net256),
    .Q(\u_rf.reg8_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12239_ (.CLK(clk),
    .D(_00276_),
    .RESET_B(net278),
    .Q(\u_rf.reg8_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12240_ (.CLK(clk),
    .D(_00277_),
    .RESET_B(net276),
    .Q(\u_rf.reg8_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12241_ (.CLK(clk),
    .D(_00278_),
    .RESET_B(net294),
    .Q(\u_rf.reg8_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12242_ (.CLK(clk),
    .D(_00279_),
    .RESET_B(net278),
    .Q(\u_rf.reg8_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12243_ (.CLK(clk),
    .D(_00280_),
    .RESET_B(net304),
    .Q(\u_rf.reg8_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12244_ (.CLK(clk),
    .D(_00281_),
    .RESET_B(net269),
    .Q(\u_rf.reg8_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12245_ (.CLK(clk),
    .D(_00282_),
    .RESET_B(net300),
    .Q(\u_rf.reg8_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12246_ (.CLK(clk),
    .D(_00283_),
    .RESET_B(net308),
    .Q(\u_rf.reg8_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12247_ (.CLK(clk),
    .D(_00284_),
    .RESET_B(net308),
    .Q(\u_rf.reg8_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12248_ (.CLK(clk),
    .D(_00285_),
    .RESET_B(net302),
    .Q(\u_rf.reg8_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12249_ (.CLK(clk),
    .D(_00286_),
    .RESET_B(net343),
    .Q(\u_rf.reg8_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12250_ (.CLK(clk),
    .D(_00287_),
    .RESET_B(net340),
    .Q(\u_rf.reg8_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12251_ (.CLK(clk),
    .D(_00288_),
    .RESET_B(net241),
    .Q(\u_rf.reg9_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12252_ (.CLK(clk),
    .D(_00289_),
    .RESET_B(net234),
    .Q(\u_rf.reg9_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12253_ (.CLK(clk),
    .D(_00290_),
    .RESET_B(net248),
    .Q(\u_rf.reg9_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12254_ (.CLK(clk),
    .D(_00291_),
    .RESET_B(net231),
    .Q(\u_rf.reg9_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12255_ (.CLK(clk),
    .D(_00292_),
    .RESET_B(net227),
    .Q(\u_rf.reg9_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12256_ (.CLK(clk),
    .D(_00293_),
    .RESET_B(net248),
    .Q(\u_rf.reg9_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12257_ (.CLK(clk),
    .D(_00294_),
    .RESET_B(net251),
    .Q(\u_rf.reg9_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12258_ (.CLK(clk),
    .D(_00295_),
    .RESET_B(net234),
    .Q(\u_rf.reg9_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12259_ (.CLK(clk),
    .D(_00296_),
    .RESET_B(net312),
    .Q(\u_rf.reg9_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12260_ (.CLK(clk),
    .D(_00297_),
    .RESET_B(net312),
    .Q(\u_rf.reg9_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12261_ (.CLK(clk),
    .D(_00298_),
    .RESET_B(net239),
    .Q(\u_rf.reg9_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12262_ (.CLK(clk),
    .D(_00299_),
    .RESET_B(net202),
    .Q(\u_rf.reg9_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12263_ (.CLK(clk),
    .D(_00300_),
    .RESET_B(net212),
    .Q(\u_rf.reg9_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12264_ (.CLK(clk),
    .D(_00301_),
    .RESET_B(net288),
    .Q(\u_rf.reg9_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12265_ (.CLK(clk),
    .D(_00302_),
    .RESET_B(net280),
    .Q(\u_rf.reg9_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12266_ (.CLK(clk),
    .D(_00303_),
    .RESET_B(net257),
    .Q(\u_rf.reg9_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12267_ (.CLK(clk),
    .D(_00304_),
    .RESET_B(net209),
    .Q(\u_rf.reg9_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12268_ (.CLK(clk),
    .D(_00305_),
    .RESET_B(net244),
    .Q(\u_rf.reg9_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12269_ (.CLK(clk),
    .D(_00306_),
    .RESET_B(net215),
    .Q(\u_rf.reg9_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12270_ (.CLK(clk),
    .D(_00307_),
    .RESET_B(net256),
    .Q(\u_rf.reg9_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12271_ (.CLK(clk),
    .D(_00308_),
    .RESET_B(net275),
    .Q(\u_rf.reg9_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12272_ (.CLK(clk),
    .D(_00309_),
    .RESET_B(net275),
    .Q(\u_rf.reg9_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12273_ (.CLK(clk),
    .D(_00310_),
    .RESET_B(net287),
    .Q(\u_rf.reg9_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12274_ (.CLK(clk),
    .D(_00311_),
    .RESET_B(net278),
    .Q(\u_rf.reg9_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12275_ (.CLK(clk),
    .D(_00312_),
    .RESET_B(net302),
    .Q(\u_rf.reg9_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12276_ (.CLK(clk),
    .D(_00313_),
    .RESET_B(net267),
    .Q(\u_rf.reg9_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12277_ (.CLK(clk),
    .D(_00314_),
    .RESET_B(net294),
    .Q(\u_rf.reg9_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12278_ (.CLK(clk),
    .D(_00315_),
    .RESET_B(net308),
    .Q(\u_rf.reg9_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12279_ (.CLK(clk),
    .D(_00316_),
    .RESET_B(net354),
    .Q(\u_rf.reg9_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12280_ (.CLK(clk),
    .D(_00317_),
    .RESET_B(net302),
    .Q(\u_rf.reg9_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12281_ (.CLK(clk),
    .D(_00318_),
    .RESET_B(net341),
    .Q(\u_rf.reg9_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12282_ (.CLK(clk),
    .D(_00319_),
    .RESET_B(net339),
    .Q(\u_rf.reg9_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12283_ (.CLK(clk),
    .D(_00320_),
    .RESET_B(net243),
    .Q(\u_rf.reg10_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12284_ (.CLK(clk),
    .D(_00321_),
    .RESET_B(net237),
    .Q(\u_rf.reg10_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12285_ (.CLK(clk),
    .D(_00322_),
    .RESET_B(net246),
    .Q(\u_rf.reg10_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12286_ (.CLK(clk),
    .D(_00323_),
    .RESET_B(net231),
    .Q(\u_rf.reg10_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12287_ (.CLK(clk),
    .D(_00324_),
    .RESET_B(net227),
    .Q(\u_rf.reg10_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12288_ (.CLK(clk),
    .D(_00325_),
    .RESET_B(net323),
    .Q(\u_rf.reg10_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12289_ (.CLK(clk),
    .D(_00326_),
    .RESET_B(net251),
    .Q(\u_rf.reg10_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12290_ (.CLK(clk),
    .D(_00327_),
    .RESET_B(net234),
    .Q(\u_rf.reg10_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12291_ (.CLK(clk),
    .D(_00328_),
    .RESET_B(net314),
    .Q(\u_rf.reg10_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12292_ (.CLK(clk),
    .D(_00329_),
    .RESET_B(net314),
    .Q(\u_rf.reg10_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12293_ (.CLK(clk),
    .D(_00330_),
    .RESET_B(net248),
    .Q(\u_rf.reg10_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12294_ (.CLK(clk),
    .D(_00331_),
    .RESET_B(net202),
    .Q(\u_rf.reg10_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12295_ (.CLK(clk),
    .D(_00332_),
    .RESET_B(net212),
    .Q(\u_rf.reg10_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12296_ (.CLK(clk),
    .D(_00333_),
    .RESET_B(net282),
    .Q(\u_rf.reg10_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12297_ (.CLK(clk),
    .D(_00334_),
    .RESET_B(net267),
    .Q(\u_rf.reg10_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12298_ (.CLK(clk),
    .D(_00335_),
    .RESET_B(net261),
    .Q(\u_rf.reg10_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12299_ (.CLK(clk),
    .D(_00336_),
    .RESET_B(net209),
    .Q(\u_rf.reg10_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12300_ (.CLK(clk),
    .D(_00337_),
    .RESET_B(net266),
    .Q(\u_rf.reg10_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12301_ (.CLK(clk),
    .D(_00338_),
    .RESET_B(net216),
    .Q(\u_rf.reg10_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12302_ (.CLK(clk),
    .D(_00339_),
    .RESET_B(net216),
    .Q(\u_rf.reg10_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12303_ (.CLK(clk),
    .D(_00340_),
    .RESET_B(net295),
    .Q(\u_rf.reg10_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12304_ (.CLK(clk),
    .D(_00341_),
    .RESET_B(net268),
    .Q(\u_rf.reg10_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12305_ (.CLK(clk),
    .D(_00342_),
    .RESET_B(net286),
    .Q(\u_rf.reg10_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12306_ (.CLK(clk),
    .D(_00343_),
    .RESET_B(net278),
    .Q(\u_rf.reg10_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12307_ (.CLK(clk),
    .D(_00344_),
    .RESET_B(net303),
    .Q(\u_rf.reg10_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12308_ (.CLK(clk),
    .D(_00345_),
    .RESET_B(net267),
    .Q(\u_rf.reg10_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12309_ (.CLK(clk),
    .D(_00346_),
    .RESET_B(net296),
    .Q(\u_rf.reg10_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12310_ (.CLK(clk),
    .D(_00347_),
    .RESET_B(net308),
    .Q(\u_rf.reg10_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12311_ (.CLK(clk),
    .D(_00348_),
    .RESET_B(net353),
    .Q(\u_rf.reg10_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12312_ (.CLK(clk),
    .D(_00349_),
    .RESET_B(net304),
    .Q(\u_rf.reg10_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12313_ (.CLK(clk),
    .D(_00350_),
    .RESET_B(net342),
    .Q(\u_rf.reg10_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12314_ (.CLK(clk),
    .D(_00351_),
    .RESET_B(net339),
    .Q(\u_rf.reg10_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12315_ (.CLK(clk),
    .D(_00352_),
    .RESET_B(net242),
    .Q(\u_rf.reg11_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12316_ (.CLK(clk),
    .D(_00353_),
    .RESET_B(net236),
    .Q(\u_rf.reg11_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12317_ (.CLK(clk),
    .D(_00354_),
    .RESET_B(net250),
    .Q(\u_rf.reg11_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12318_ (.CLK(clk),
    .D(_00355_),
    .RESET_B(net241),
    .Q(\u_rf.reg11_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12319_ (.CLK(clk),
    .D(_00356_),
    .RESET_B(net227),
    .Q(\u_rf.reg11_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12320_ (.CLK(clk),
    .D(_00357_),
    .RESET_B(net323),
    .Q(\u_rf.reg11_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12321_ (.CLK(clk),
    .D(_00358_),
    .RESET_B(net326),
    .Q(\u_rf.reg11_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12322_ (.CLK(clk),
    .D(_00359_),
    .RESET_B(net234),
    .Q(\u_rf.reg11_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12323_ (.CLK(clk),
    .D(_00360_),
    .RESET_B(net313),
    .Q(\u_rf.reg11_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12324_ (.CLK(clk),
    .D(_00361_),
    .RESET_B(net313),
    .Q(\u_rf.reg11_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12325_ (.CLK(clk),
    .D(_00362_),
    .RESET_B(net240),
    .Q(\u_rf.reg11_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12326_ (.CLK(clk),
    .D(_00363_),
    .RESET_B(net210),
    .Q(\u_rf.reg11_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12327_ (.CLK(clk),
    .D(_00364_),
    .RESET_B(net213),
    .Q(\u_rf.reg11_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12328_ (.CLK(clk),
    .D(_00365_),
    .RESET_B(net291),
    .Q(\u_rf.reg11_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12329_ (.CLK(clk),
    .D(_00366_),
    .RESET_B(net286),
    .Q(\u_rf.reg11_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12330_ (.CLK(clk),
    .D(_00367_),
    .RESET_B(net262),
    .Q(\u_rf.reg11_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12331_ (.CLK(clk),
    .D(_00368_),
    .RESET_B(net205),
    .Q(\u_rf.reg11_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12332_ (.CLK(clk),
    .D(_00369_),
    .RESET_B(net246),
    .Q(\u_rf.reg11_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12333_ (.CLK(clk),
    .D(_00370_),
    .RESET_B(net217),
    .Q(\u_rf.reg11_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12334_ (.CLK(clk),
    .D(_00371_),
    .RESET_B(net258),
    .Q(\u_rf.reg11_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12335_ (.CLK(clk),
    .D(_00372_),
    .RESET_B(net294),
    .Q(\u_rf.reg11_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12336_ (.CLK(clk),
    .D(_00373_),
    .RESET_B(net275),
    .Q(\u_rf.reg11_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12337_ (.CLK(clk),
    .D(_00374_),
    .RESET_B(net285),
    .Q(\u_rf.reg11_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12338_ (.CLK(clk),
    .D(_00375_),
    .RESET_B(net298),
    .Q(\u_rf.reg11_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12339_ (.CLK(clk),
    .D(_00376_),
    .RESET_B(net304),
    .Q(\u_rf.reg11_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12340_ (.CLK(clk),
    .D(_00377_),
    .RESET_B(net268),
    .Q(\u_rf.reg11_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12341_ (.CLK(clk),
    .D(_00378_),
    .RESET_B(net298),
    .Q(\u_rf.reg11_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12342_ (.CLK(clk),
    .D(_00379_),
    .RESET_B(net308),
    .Q(\u_rf.reg11_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12343_ (.CLK(clk),
    .D(_00380_),
    .RESET_B(net352),
    .Q(\u_rf.reg11_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12344_ (.CLK(clk),
    .D(_00381_),
    .RESET_B(net342),
    .Q(\u_rf.reg11_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12345_ (.CLK(clk),
    .D(_00382_),
    .RESET_B(net293),
    .Q(\u_rf.reg11_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12346_ (.CLK(clk),
    .D(_00383_),
    .RESET_B(net341),
    .Q(\u_rf.reg11_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12347_ (.CLK(clk),
    .D(_00384_),
    .RESET_B(net243),
    .Q(\u_rf.reg12_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12348_ (.CLK(clk),
    .D(_00385_),
    .RESET_B(net237),
    .Q(\u_rf.reg12_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12349_ (.CLK(clk),
    .D(_00386_),
    .RESET_B(net245),
    .Q(\u_rf.reg12_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12350_ (.CLK(clk),
    .D(_00387_),
    .RESET_B(net231),
    .Q(\u_rf.reg12_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12351_ (.CLK(clk),
    .D(_00388_),
    .RESET_B(net228),
    .Q(\u_rf.reg12_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12352_ (.CLK(clk),
    .D(_00389_),
    .RESET_B(net323),
    .Q(\u_rf.reg12_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12353_ (.CLK(clk),
    .D(_00390_),
    .RESET_B(net251),
    .Q(\u_rf.reg12_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12354_ (.CLK(clk),
    .D(_00391_),
    .RESET_B(net229),
    .Q(\u_rf.reg12_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12355_ (.CLK(clk),
    .D(_00392_),
    .RESET_B(net314),
    .Q(\u_rf.reg12_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12356_ (.CLK(clk),
    .D(_00393_),
    .RESET_B(net317),
    .Q(\u_rf.reg12_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12357_ (.CLK(clk),
    .D(_00394_),
    .RESET_B(net248),
    .Q(\u_rf.reg12_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12358_ (.CLK(clk),
    .D(_00395_),
    .RESET_B(net204),
    .Q(\u_rf.reg12_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12359_ (.CLK(clk),
    .D(_00396_),
    .RESET_B(net212),
    .Q(\u_rf.reg12_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12360_ (.CLK(clk),
    .D(_00397_),
    .RESET_B(net289),
    .Q(\u_rf.reg12_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12361_ (.CLK(clk),
    .D(_00398_),
    .RESET_B(net280),
    .Q(\u_rf.reg12_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12362_ (.CLK(clk),
    .D(_00399_),
    .RESET_B(net257),
    .Q(\u_rf.reg12_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12363_ (.CLK(clk),
    .D(_00400_),
    .RESET_B(net208),
    .Q(\u_rf.reg12_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12364_ (.CLK(clk),
    .D(_00401_),
    .RESET_B(net280),
    .Q(\u_rf.reg12_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12365_ (.CLK(clk),
    .D(_00402_),
    .RESET_B(net215),
    .Q(\u_rf.reg12_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12366_ (.CLK(clk),
    .D(_00403_),
    .RESET_B(net216),
    .Q(\u_rf.reg12_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12367_ (.CLK(clk),
    .D(_00404_),
    .RESET_B(net276),
    .Q(\u_rf.reg12_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12368_ (.CLK(clk),
    .D(_00405_),
    .RESET_B(net276),
    .Q(\u_rf.reg12_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12369_ (.CLK(clk),
    .D(_00406_),
    .RESET_B(net287),
    .Q(\u_rf.reg12_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12370_ (.CLK(clk),
    .D(_00407_),
    .RESET_B(net277),
    .Q(\u_rf.reg12_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12371_ (.CLK(clk),
    .D(_00408_),
    .RESET_B(net350),
    .Q(\u_rf.reg12_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12372_ (.CLK(clk),
    .D(_00409_),
    .RESET_B(net269),
    .Q(\u_rf.reg12_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12373_ (.CLK(clk),
    .D(_00410_),
    .RESET_B(net296),
    .Q(\u_rf.reg12_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12374_ (.CLK(clk),
    .D(_00411_),
    .RESET_B(net307),
    .Q(\u_rf.reg12_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12375_ (.CLK(clk),
    .D(_00412_),
    .RESET_B(net353),
    .Q(\u_rf.reg12_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12376_ (.CLK(clk),
    .D(_00413_),
    .RESET_B(net342),
    .Q(\u_rf.reg12_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12377_ (.CLK(clk),
    .D(_00414_),
    .RESET_B(net292),
    .Q(\u_rf.reg12_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12378_ (.CLK(clk),
    .D(_00415_),
    .RESET_B(net340),
    .Q(\u_rf.reg12_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12379_ (.CLK(clk),
    .D(_00416_),
    .RESET_B(net222),
    .Q(\u_rf.reg13_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12380_ (.CLK(clk),
    .D(_00417_),
    .RESET_B(net240),
    .Q(\u_rf.reg13_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12381_ (.CLK(clk),
    .D(_00418_),
    .RESET_B(net245),
    .Q(\u_rf.reg13_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12382_ (.CLK(clk),
    .D(_00419_),
    .RESET_B(net232),
    .Q(\u_rf.reg13_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12383_ (.CLK(clk),
    .D(_00420_),
    .RESET_B(net205),
    .Q(\u_rf.reg13_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12384_ (.CLK(clk),
    .D(_00421_),
    .RESET_B(net323),
    .Q(\u_rf.reg13_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12385_ (.CLK(clk),
    .D(_00422_),
    .RESET_B(net325),
    .Q(\u_rf.reg13_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12386_ (.CLK(clk),
    .D(_00423_),
    .RESET_B(net229),
    .Q(\u_rf.reg13_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12387_ (.CLK(clk),
    .D(_00424_),
    .RESET_B(net315),
    .Q(\u_rf.reg13_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12388_ (.CLK(clk),
    .D(_00425_),
    .RESET_B(net317),
    .Q(\u_rf.reg13_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12389_ (.CLK(clk),
    .D(_00426_),
    .RESET_B(net241),
    .Q(\u_rf.reg13_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12390_ (.CLK(clk),
    .D(_00427_),
    .RESET_B(net203),
    .Q(\u_rf.reg13_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12391_ (.CLK(clk),
    .D(_00428_),
    .RESET_B(net213),
    .Q(\u_rf.reg13_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12392_ (.CLK(clk),
    .D(_00429_),
    .RESET_B(net291),
    .Q(\u_rf.reg13_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12393_ (.CLK(clk),
    .D(_00430_),
    .RESET_B(net286),
    .Q(\u_rf.reg13_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12394_ (.CLK(clk),
    .D(_00431_),
    .RESET_B(net269),
    .Q(\u_rf.reg13_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12395_ (.CLK(clk),
    .D(_00432_),
    .RESET_B(net207),
    .Q(\u_rf.reg13_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12396_ (.CLK(clk),
    .D(_00433_),
    .RESET_B(net225),
    .Q(\u_rf.reg13_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12397_ (.CLK(clk),
    .D(_00434_),
    .RESET_B(net217),
    .Q(\u_rf.reg13_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12398_ (.CLK(clk),
    .D(_00435_),
    .RESET_B(net258),
    .Q(\u_rf.reg13_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12399_ (.CLK(clk),
    .D(_00436_),
    .RESET_B(net273),
    .Q(\u_rf.reg13_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12400_ (.CLK(clk),
    .D(_00437_),
    .RESET_B(net273),
    .Q(\u_rf.reg13_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12401_ (.CLK(clk),
    .D(_00438_),
    .RESET_B(net302),
    .Q(\u_rf.reg13_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12402_ (.CLK(clk),
    .D(_00439_),
    .RESET_B(net278),
    .Q(\u_rf.reg13_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12403_ (.CLK(clk),
    .D(_00440_),
    .RESET_B(net302),
    .Q(\u_rf.reg13_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12404_ (.CLK(clk),
    .D(_00441_),
    .RESET_B(net261),
    .Q(\u_rf.reg13_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12405_ (.CLK(clk),
    .D(_00442_),
    .RESET_B(net298),
    .Q(\u_rf.reg13_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12406_ (.CLK(clk),
    .D(_00443_),
    .RESET_B(net306),
    .Q(\u_rf.reg13_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12407_ (.CLK(clk),
    .D(_00444_),
    .RESET_B(net352),
    .Q(\u_rf.reg13_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12408_ (.CLK(clk),
    .D(_00445_),
    .RESET_B(net304),
    .Q(\u_rf.reg13_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12409_ (.CLK(clk),
    .D(_00446_),
    .RESET_B(net343),
    .Q(\u_rf.reg13_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12410_ (.CLK(clk),
    .D(_00447_),
    .RESET_B(net343),
    .Q(\u_rf.reg13_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12411_ (.CLK(clk),
    .D(_00448_),
    .RESET_B(net243),
    .Q(\u_rf.reg14_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12412_ (.CLK(clk),
    .D(_00449_),
    .RESET_B(net236),
    .Q(\u_rf.reg14_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12413_ (.CLK(clk),
    .D(_00450_),
    .RESET_B(net245),
    .Q(\u_rf.reg14_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12414_ (.CLK(clk),
    .D(_00451_),
    .RESET_B(net243),
    .Q(\u_rf.reg14_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12415_ (.CLK(clk),
    .D(_00452_),
    .RESET_B(net227),
    .Q(\u_rf.reg14_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12416_ (.CLK(clk),
    .D(_00453_),
    .RESET_B(net248),
    .Q(\u_rf.reg14_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12417_ (.CLK(clk),
    .D(_00454_),
    .RESET_B(net251),
    .Q(\u_rf.reg14_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12418_ (.CLK(clk),
    .D(_00455_),
    .RESET_B(net230),
    .Q(\u_rf.reg14_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12419_ (.CLK(clk),
    .D(_00456_),
    .RESET_B(net312),
    .Q(\u_rf.reg14_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12420_ (.CLK(clk),
    .D(_00457_),
    .RESET_B(net313),
    .Q(\u_rf.reg14_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12421_ (.CLK(clk),
    .D(_00458_),
    .RESET_B(net241),
    .Q(\u_rf.reg14_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12422_ (.CLK(clk),
    .D(_00459_),
    .RESET_B(net203),
    .Q(\u_rf.reg14_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12423_ (.CLK(clk),
    .D(_00460_),
    .RESET_B(net213),
    .Q(\u_rf.reg14_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12424_ (.CLK(clk),
    .D(_00461_),
    .RESET_B(net289),
    .Q(\u_rf.reg14_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12425_ (.CLK(clk),
    .D(_00462_),
    .RESET_B(net282),
    .Q(\u_rf.reg14_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12426_ (.CLK(clk),
    .D(_00463_),
    .RESET_B(net258),
    .Q(\u_rf.reg14_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12427_ (.CLK(clk),
    .D(_00464_),
    .RESET_B(net221),
    .Q(\u_rf.reg14_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12428_ (.CLK(clk),
    .D(_00465_),
    .RESET_B(net281),
    .Q(\u_rf.reg14_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12429_ (.CLK(clk),
    .D(_00466_),
    .RESET_B(net217),
    .Q(\u_rf.reg14_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12430_ (.CLK(clk),
    .D(_00467_),
    .RESET_B(net258),
    .Q(\u_rf.reg14_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12431_ (.CLK(clk),
    .D(_00468_),
    .RESET_B(net273),
    .Q(\u_rf.reg14_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12432_ (.CLK(clk),
    .D(_00469_),
    .RESET_B(net273),
    .Q(\u_rf.reg14_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12433_ (.CLK(clk),
    .D(_00470_),
    .RESET_B(net302),
    .Q(\u_rf.reg14_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12434_ (.CLK(clk),
    .D(_00471_),
    .RESET_B(net277),
    .Q(\u_rf.reg14_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12435_ (.CLK(clk),
    .D(_00472_),
    .RESET_B(net350),
    .Q(\u_rf.reg14_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12436_ (.CLK(clk),
    .D(_00473_),
    .RESET_B(net261),
    .Q(\u_rf.reg14_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12437_ (.CLK(clk),
    .D(_00474_),
    .RESET_B(net300),
    .Q(\u_rf.reg14_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12438_ (.CLK(clk),
    .D(_00475_),
    .RESET_B(net306),
    .Q(\u_rf.reg14_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12439_ (.CLK(clk),
    .D(_00476_),
    .RESET_B(net353),
    .Q(\u_rf.reg14_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12440_ (.CLK(clk),
    .D(_00477_),
    .RESET_B(net349),
    .Q(\u_rf.reg14_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12441_ (.CLK(clk),
    .D(_00478_),
    .RESET_B(net292),
    .Q(\u_rf.reg14_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12442_ (.CLK(clk),
    .D(_00479_),
    .RESET_B(net340),
    .Q(\u_rf.reg14_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12443_ (.CLK(clk),
    .D(_00480_),
    .RESET_B(net222),
    .Q(\u_rf.reg15_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12444_ (.CLK(clk),
    .D(_00481_),
    .RESET_B(net236),
    .Q(\u_rf.reg15_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12445_ (.CLK(clk),
    .D(_00482_),
    .RESET_B(net245),
    .Q(\u_rf.reg15_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12446_ (.CLK(clk),
    .D(_00483_),
    .RESET_B(net205),
    .Q(\u_rf.reg15_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12447_ (.CLK(clk),
    .D(_00484_),
    .RESET_B(net206),
    .Q(\u_rf.reg15_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12448_ (.CLK(clk),
    .D(_00485_),
    .RESET_B(net324),
    .Q(\u_rf.reg15_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12449_ (.CLK(clk),
    .D(_00486_),
    .RESET_B(net326),
    .Q(\u_rf.reg15_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12450_ (.CLK(clk),
    .D(_00487_),
    .RESET_B(net229),
    .Q(\u_rf.reg15_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12451_ (.CLK(clk),
    .D(_00488_),
    .RESET_B(net312),
    .Q(\u_rf.reg15_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12452_ (.CLK(clk),
    .D(_00489_),
    .RESET_B(net316),
    .Q(\u_rf.reg15_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12453_ (.CLK(clk),
    .D(_00490_),
    .RESET_B(net247),
    .Q(\u_rf.reg15_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12454_ (.CLK(clk),
    .D(_00491_),
    .RESET_B(net210),
    .Q(\u_rf.reg15_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12455_ (.CLK(clk),
    .D(_00492_),
    .RESET_B(net223),
    .Q(\u_rf.reg15_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12456_ (.CLK(clk),
    .D(_00493_),
    .RESET_B(net288),
    .Q(\u_rf.reg15_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12457_ (.CLK(clk),
    .D(_00494_),
    .RESET_B(net286),
    .Q(\u_rf.reg15_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12458_ (.CLK(clk),
    .D(_00495_),
    .RESET_B(net266),
    .Q(\u_rf.reg15_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12459_ (.CLK(clk),
    .D(_00496_),
    .RESET_B(net207),
    .Q(\u_rf.reg15_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12460_ (.CLK(clk),
    .D(_00497_),
    .RESET_B(net280),
    .Q(\u_rf.reg15_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12461_ (.CLK(clk),
    .D(_00498_),
    .RESET_B(net226),
    .Q(\u_rf.reg15_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12462_ (.CLK(clk),
    .D(_00499_),
    .RESET_B(net258),
    .Q(\u_rf.reg15_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12463_ (.CLK(clk),
    .D(_00500_),
    .RESET_B(net273),
    .Q(\u_rf.reg15_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12464_ (.CLK(clk),
    .D(_00501_),
    .RESET_B(net273),
    .Q(\u_rf.reg15_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12465_ (.CLK(clk),
    .D(_00502_),
    .RESET_B(net296),
    .Q(\u_rf.reg15_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12466_ (.CLK(clk),
    .D(_00503_),
    .RESET_B(net277),
    .Q(\u_rf.reg15_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12467_ (.CLK(clk),
    .D(_00504_),
    .RESET_B(net305),
    .Q(\u_rf.reg15_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12468_ (.CLK(clk),
    .D(_00505_),
    .RESET_B(net261),
    .Q(\u_rf.reg15_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12469_ (.CLK(clk),
    .D(_00506_),
    .RESET_B(net300),
    .Q(\u_rf.reg15_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12470_ (.CLK(clk),
    .D(_00507_),
    .RESET_B(net306),
    .Q(\u_rf.reg15_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12471_ (.CLK(clk),
    .D(_00508_),
    .RESET_B(net353),
    .Q(\u_rf.reg15_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12472_ (.CLK(clk),
    .D(_00509_),
    .RESET_B(net349),
    .Q(\u_rf.reg15_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12473_ (.CLK(clk),
    .D(_00510_),
    .RESET_B(net293),
    .Q(\u_rf.reg15_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12474_ (.CLK(clk),
    .D(_00511_),
    .RESET_B(net339),
    .Q(\u_rf.reg15_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12475_ (.CLK(clk),
    .D(_00512_),
    .RESET_B(net224),
    .Q(\u_rf.reg16_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12476_ (.CLK(clk),
    .D(_00513_),
    .RESET_B(net237),
    .Q(\u_rf.reg16_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12477_ (.CLK(clk),
    .D(_00514_),
    .RESET_B(net244),
    .Q(\u_rf.reg16_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12478_ (.CLK(clk),
    .D(_00515_),
    .RESET_B(net232),
    .Q(\u_rf.reg16_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12479_ (.CLK(clk),
    .D(_00516_),
    .RESET_B(net205),
    .Q(\u_rf.reg16_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12480_ (.CLK(clk),
    .D(_00517_),
    .RESET_B(net324),
    .Q(\u_rf.reg16_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12481_ (.CLK(clk),
    .D(_00518_),
    .RESET_B(net326),
    .Q(\u_rf.reg16_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12482_ (.CLK(clk),
    .D(_00519_),
    .RESET_B(net230),
    .Q(\u_rf.reg16_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12483_ (.CLK(clk),
    .D(_00520_),
    .RESET_B(net313),
    .Q(\u_rf.reg16_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12484_ (.CLK(clk),
    .D(_00521_),
    .RESET_B(net316),
    .Q(\u_rf.reg16_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12485_ (.CLK(clk),
    .D(_00522_),
    .RESET_B(net239),
    .Q(\u_rf.reg16_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12486_ (.CLK(clk),
    .D(_00523_),
    .RESET_B(net203),
    .Q(\u_rf.reg16_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12487_ (.CLK(clk),
    .D(_00524_),
    .RESET_B(net213),
    .Q(\u_rf.reg16_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12488_ (.CLK(clk),
    .D(_00525_),
    .RESET_B(net289),
    .Q(\u_rf.reg16_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12489_ (.CLK(clk),
    .D(_00526_),
    .RESET_B(net270),
    .Q(\u_rf.reg16_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12490_ (.CLK(clk),
    .D(_00527_),
    .RESET_B(net259),
    .Q(\u_rf.reg16_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12491_ (.CLK(clk),
    .D(_00528_),
    .RESET_B(net208),
    .Q(\u_rf.reg16_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12492_ (.CLK(clk),
    .D(_00529_),
    .RESET_B(net265),
    .Q(\u_rf.reg16_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12493_ (.CLK(clk),
    .D(_00530_),
    .RESET_B(net217),
    .Q(\u_rf.reg16_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12494_ (.CLK(clk),
    .D(_00531_),
    .RESET_B(net218),
    .Q(\u_rf.reg16_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12495_ (.CLK(clk),
    .D(_00532_),
    .RESET_B(net274),
    .Q(\u_rf.reg16_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12496_ (.CLK(clk),
    .D(_00533_),
    .RESET_B(net263),
    .Q(\u_rf.reg16_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12497_ (.CLK(clk),
    .D(_00534_),
    .RESET_B(net302),
    .Q(\u_rf.reg16_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12498_ (.CLK(clk),
    .D(_00535_),
    .RESET_B(net274),
    .Q(\u_rf.reg16_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12499_ (.CLK(clk),
    .D(_00536_),
    .RESET_B(net350),
    .Q(\u_rf.reg16_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12500_ (.CLK(clk),
    .D(_00537_),
    .RESET_B(net263),
    .Q(\u_rf.reg16_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12501_ (.CLK(clk),
    .D(_00538_),
    .RESET_B(net298),
    .Q(\u_rf.reg16_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12502_ (.CLK(clk),
    .D(_00539_),
    .RESET_B(net300),
    .Q(\u_rf.reg16_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12503_ (.CLK(clk),
    .D(_00540_),
    .RESET_B(net352),
    .Q(\u_rf.reg16_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12504_ (.CLK(clk),
    .D(_00541_),
    .RESET_B(net304),
    .Q(\u_rf.reg16_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12505_ (.CLK(clk),
    .D(_00542_),
    .RESET_B(net292),
    .Q(\u_rf.reg16_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12506_ (.CLK(clk),
    .D(_00543_),
    .RESET_B(net292),
    .Q(\u_rf.reg16_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12507_ (.CLK(clk),
    .D(_00544_),
    .RESET_B(net221),
    .Q(\u_rf.reg17_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12508_ (.CLK(clk),
    .D(_00545_),
    .RESET_B(net237),
    .Q(\u_rf.reg17_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12509_ (.CLK(clk),
    .D(_00546_),
    .RESET_B(net224),
    .Q(\u_rf.reg17_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12510_ (.CLK(clk),
    .D(_00547_),
    .RESET_B(net209),
    .Q(\u_rf.reg17_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12511_ (.CLK(clk),
    .D(_00548_),
    .RESET_B(net205),
    .Q(\u_rf.reg17_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12512_ (.CLK(clk),
    .D(_00549_),
    .RESET_B(net323),
    .Q(\u_rf.reg17_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12513_ (.CLK(clk),
    .D(_00550_),
    .RESET_B(net251),
    .Q(\u_rf.reg17_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12514_ (.CLK(clk),
    .D(_00551_),
    .RESET_B(net231),
    .Q(\u_rf.reg17_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12515_ (.CLK(clk),
    .D(_00552_),
    .RESET_B(net315),
    .Q(\u_rf.reg17_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12516_ (.CLK(clk),
    .D(_00553_),
    .RESET_B(net317),
    .Q(\u_rf.reg17_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12517_ (.CLK(clk),
    .D(_00554_),
    .RESET_B(net239),
    .Q(\u_rf.reg17_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12518_ (.CLK(clk),
    .D(_00555_),
    .RESET_B(net203),
    .Q(\u_rf.reg17_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12519_ (.CLK(clk),
    .D(_00556_),
    .RESET_B(net212),
    .Q(\u_rf.reg17_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12520_ (.CLK(clk),
    .D(_00557_),
    .RESET_B(net288),
    .Q(\u_rf.reg17_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12521_ (.CLK(clk),
    .D(_00558_),
    .RESET_B(net267),
    .Q(\u_rf.reg17_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12522_ (.CLK(clk),
    .D(_00559_),
    .RESET_B(net261),
    .Q(\u_rf.reg17_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12523_ (.CLK(clk),
    .D(_00560_),
    .RESET_B(net205),
    .Q(\u_rf.reg17_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12524_ (.CLK(clk),
    .D(_00561_),
    .RESET_B(net225),
    .Q(\u_rf.reg17_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12525_ (.CLK(clk),
    .D(_00562_),
    .RESET_B(net216),
    .Q(\u_rf.reg17_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12526_ (.CLK(clk),
    .D(_00563_),
    .RESET_B(net256),
    .Q(\u_rf.reg17_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12527_ (.CLK(clk),
    .D(_00564_),
    .RESET_B(net274),
    .Q(\u_rf.reg17_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12528_ (.CLK(clk),
    .D(_00565_),
    .RESET_B(net263),
    .Q(\u_rf.reg17_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12529_ (.CLK(clk),
    .D(_00566_),
    .RESET_B(net296),
    .Q(\u_rf.reg17_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12530_ (.CLK(clk),
    .D(_00567_),
    .RESET_B(net274),
    .Q(\u_rf.reg17_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12531_ (.CLK(clk),
    .D(_00568_),
    .RESET_B(net305),
    .Q(\u_rf.reg17_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12532_ (.CLK(clk),
    .D(_00569_),
    .RESET_B(net262),
    .Q(\u_rf.reg17_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12533_ (.CLK(clk),
    .D(_00570_),
    .RESET_B(net295),
    .Q(\u_rf.reg17_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12534_ (.CLK(clk),
    .D(_00571_),
    .RESET_B(net300),
    .Q(\u_rf.reg17_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12535_ (.CLK(clk),
    .D(_00572_),
    .RESET_B(net353),
    .Q(\u_rf.reg17_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12536_ (.CLK(clk),
    .D(_00573_),
    .RESET_B(net349),
    .Q(\u_rf.reg17_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12537_ (.CLK(clk),
    .D(_00574_),
    .RESET_B(net293),
    .Q(\u_rf.reg17_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12538_ (.CLK(clk),
    .D(_00575_),
    .RESET_B(net289),
    .Q(\u_rf.reg17_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12539_ (.CLK(clk),
    .D(_00576_),
    .RESET_B(net243),
    .Q(\u_rf.reg18_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12540_ (.CLK(clk),
    .D(_00577_),
    .RESET_B(net235),
    .Q(\u_rf.reg18_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12541_ (.CLK(clk),
    .D(_00578_),
    .RESET_B(net245),
    .Q(\u_rf.reg18_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12542_ (.CLK(clk),
    .D(_00579_),
    .RESET_B(net232),
    .Q(\u_rf.reg18_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12543_ (.CLK(clk),
    .D(_00580_),
    .RESET_B(net228),
    .Q(\u_rf.reg18_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12544_ (.CLK(clk),
    .D(_00581_),
    .RESET_B(net323),
    .Q(\u_rf.reg18_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12545_ (.CLK(clk),
    .D(_00582_),
    .RESET_B(net325),
    .Q(\u_rf.reg18_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12546_ (.CLK(clk),
    .D(_00583_),
    .RESET_B(net230),
    .Q(\u_rf.reg18_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12547_ (.CLK(clk),
    .D(_00584_),
    .RESET_B(net319),
    .Q(\u_rf.reg18_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12548_ (.CLK(clk),
    .D(_00585_),
    .RESET_B(net321),
    .Q(\u_rf.reg18_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12549_ (.CLK(clk),
    .D(_00586_),
    .RESET_B(net316),
    .Q(\u_rf.reg18_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12550_ (.CLK(clk),
    .D(_00587_),
    .RESET_B(net203),
    .Q(\u_rf.reg18_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12551_ (.CLK(clk),
    .D(_00588_),
    .RESET_B(net212),
    .Q(\u_rf.reg18_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12552_ (.CLK(clk),
    .D(_00589_),
    .RESET_B(net288),
    .Q(\u_rf.reg18_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12553_ (.CLK(clk),
    .D(_00590_),
    .RESET_B(net284),
    .Q(\u_rf.reg18_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12554_ (.CLK(clk),
    .D(_00591_),
    .RESET_B(net261),
    .Q(\u_rf.reg18_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12555_ (.CLK(clk),
    .D(_00592_),
    .RESET_B(net209),
    .Q(\u_rf.reg18_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12556_ (.CLK(clk),
    .D(_00593_),
    .RESET_B(net225),
    .Q(\u_rf.reg18_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12557_ (.CLK(clk),
    .D(_00594_),
    .RESET_B(net216),
    .Q(\u_rf.reg18_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12558_ (.CLK(clk),
    .D(_00595_),
    .RESET_B(net256),
    .Q(\u_rf.reg18_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12559_ (.CLK(clk),
    .D(_00596_),
    .RESET_B(net275),
    .Q(\u_rf.reg18_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12560_ (.CLK(clk),
    .D(_00597_),
    .RESET_B(net269),
    .Q(\u_rf.reg18_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12561_ (.CLK(clk),
    .D(_00598_),
    .RESET_B(net291),
    .Q(\u_rf.reg18_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12562_ (.CLK(clk),
    .D(_00599_),
    .RESET_B(net278),
    .Q(\u_rf.reg18_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12563_ (.CLK(clk),
    .D(_00600_),
    .RESET_B(net351),
    .Q(\u_rf.reg18_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12564_ (.CLK(clk),
    .D(_00601_),
    .RESET_B(net267),
    .Q(\u_rf.reg18_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12565_ (.CLK(clk),
    .D(_00602_),
    .RESET_B(net299),
    .Q(\u_rf.reg18_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12566_ (.CLK(clk),
    .D(_00603_),
    .RESET_B(net308),
    .Q(\u_rf.reg18_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12567_ (.CLK(clk),
    .D(_00604_),
    .RESET_B(net352),
    .Q(\u_rf.reg18_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12568_ (.CLK(clk),
    .D(_00605_),
    .RESET_B(net351),
    .Q(\u_rf.reg18_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12569_ (.CLK(clk),
    .D(_00606_),
    .RESET_B(net341),
    .Q(\u_rf.reg18_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12570_ (.CLK(clk),
    .D(_00607_),
    .RESET_B(net346),
    .Q(\u_rf.reg18_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12571_ (.CLK(clk),
    .D(_00608_),
    .RESET_B(net222),
    .Q(\u_rf.reg19_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12572_ (.CLK(clk),
    .D(_00609_),
    .RESET_B(net237),
    .Q(\u_rf.reg19_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12573_ (.CLK(clk),
    .D(_00610_),
    .RESET_B(net244),
    .Q(\u_rf.reg19_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12574_ (.CLK(clk),
    .D(_00611_),
    .RESET_B(net221),
    .Q(\u_rf.reg19_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12575_ (.CLK(clk),
    .D(_00612_),
    .RESET_B(net205),
    .Q(\u_rf.reg19_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12576_ (.CLK(clk),
    .D(_00613_),
    .RESET_B(net324),
    .Q(\u_rf.reg19_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12577_ (.CLK(clk),
    .D(_00614_),
    .RESET_B(net326),
    .Q(\u_rf.reg19_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12578_ (.CLK(clk),
    .D(_00615_),
    .RESET_B(net230),
    .Q(\u_rf.reg19_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12579_ (.CLK(clk),
    .D(_00616_),
    .RESET_B(net313),
    .Q(\u_rf.reg19_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12580_ (.CLK(clk),
    .D(_00617_),
    .RESET_B(net316),
    .Q(\u_rf.reg19_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12581_ (.CLK(clk),
    .D(_00618_),
    .RESET_B(net239),
    .Q(\u_rf.reg19_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12582_ (.CLK(clk),
    .D(_00619_),
    .RESET_B(net204),
    .Q(\u_rf.reg19_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12583_ (.CLK(clk),
    .D(_00620_),
    .RESET_B(net214),
    .Q(\u_rf.reg19_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12584_ (.CLK(clk),
    .D(_00621_),
    .RESET_B(net281),
    .Q(\u_rf.reg19_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12585_ (.CLK(clk),
    .D(_00622_),
    .RESET_B(net280),
    .Q(\u_rf.reg19_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12586_ (.CLK(clk),
    .D(_00623_),
    .RESET_B(net259),
    .Q(\u_rf.reg19_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12587_ (.CLK(clk),
    .D(_00624_),
    .RESET_B(net208),
    .Q(\u_rf.reg19_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12588_ (.CLK(clk),
    .D(_00625_),
    .RESET_B(net265),
    .Q(\u_rf.reg19_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12589_ (.CLK(clk),
    .D(_00626_),
    .RESET_B(net217),
    .Q(\u_rf.reg19_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12590_ (.CLK(clk),
    .D(_00627_),
    .RESET_B(net219),
    .Q(\u_rf.reg19_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12591_ (.CLK(clk),
    .D(_00628_),
    .RESET_B(net274),
    .Q(\u_rf.reg19_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12592_ (.CLK(clk),
    .D(_00629_),
    .RESET_B(net263),
    .Q(\u_rf.reg19_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12593_ (.CLK(clk),
    .D(_00630_),
    .RESET_B(net286),
    .Q(\u_rf.reg19_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12594_ (.CLK(clk),
    .D(_00631_),
    .RESET_B(net274),
    .Q(\u_rf.reg19_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12595_ (.CLK(clk),
    .D(_00632_),
    .RESET_B(net350),
    .Q(\u_rf.reg19_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12596_ (.CLK(clk),
    .D(_00633_),
    .RESET_B(net263),
    .Q(\u_rf.reg19_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12597_ (.CLK(clk),
    .D(_00634_),
    .RESET_B(net299),
    .Q(\u_rf.reg19_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12598_ (.CLK(clk),
    .D(_00635_),
    .RESET_B(net306),
    .Q(\u_rf.reg19_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12599_ (.CLK(clk),
    .D(_00636_),
    .RESET_B(net353),
    .Q(\u_rf.reg19_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12600_ (.CLK(clk),
    .D(_00637_),
    .RESET_B(net342),
    .Q(\u_rf.reg19_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12601_ (.CLK(clk),
    .D(_00638_),
    .RESET_B(net343),
    .Q(\u_rf.reg19_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12602_ (.CLK(clk),
    .D(_00639_),
    .RESET_B(net292),
    .Q(\u_rf.reg19_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12603_ (.CLK(clk),
    .D(_00640_),
    .RESET_B(net241),
    .Q(\u_rf.reg20_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12604_ (.CLK(clk),
    .D(_00641_),
    .RESET_B(net235),
    .Q(\u_rf.reg20_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12605_ (.CLK(clk),
    .D(_00642_),
    .RESET_B(net246),
    .Q(\u_rf.reg20_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12606_ (.CLK(clk),
    .D(_00643_),
    .RESET_B(net231),
    .Q(\u_rf.reg20_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12607_ (.CLK(clk),
    .D(_00644_),
    .RESET_B(net228),
    .Q(\u_rf.reg20_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12608_ (.CLK(clk),
    .D(_00645_),
    .RESET_B(net324),
    .Q(\u_rf.reg20_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12609_ (.CLK(clk),
    .D(_00646_),
    .RESET_B(net326),
    .Q(\u_rf.reg20_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12610_ (.CLK(clk),
    .D(_00647_),
    .RESET_B(net235),
    .Q(\u_rf.reg20_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12611_ (.CLK(clk),
    .D(_00648_),
    .RESET_B(net313),
    .Q(\u_rf.reg20_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12612_ (.CLK(clk),
    .D(_00649_),
    .RESET_B(net316),
    .Q(\u_rf.reg20_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12613_ (.CLK(clk),
    .D(_00650_),
    .RESET_B(net316),
    .Q(\u_rf.reg20_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12614_ (.CLK(clk),
    .D(_00651_),
    .RESET_B(net203),
    .Q(\u_rf.reg20_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12615_ (.CLK(clk),
    .D(_00652_),
    .RESET_B(net214),
    .Q(\u_rf.reg20_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12616_ (.CLK(clk),
    .D(_00653_),
    .RESET_B(net282),
    .Q(\u_rf.reg20_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12617_ (.CLK(clk),
    .D(_00654_),
    .RESET_B(net284),
    .Q(\u_rf.reg20_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12618_ (.CLK(clk),
    .D(_00655_),
    .RESET_B(net262),
    .Q(\u_rf.reg20_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12619_ (.CLK(clk),
    .D(_00656_),
    .RESET_B(net208),
    .Q(\u_rf.reg20_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12620_ (.CLK(clk),
    .D(_00657_),
    .RESET_B(net225),
    .Q(\u_rf.reg20_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12621_ (.CLK(clk),
    .D(_00658_),
    .RESET_B(net217),
    .Q(\u_rf.reg20_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12622_ (.CLK(clk),
    .D(_00659_),
    .RESET_B(net258),
    .Q(\u_rf.reg20_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12623_ (.CLK(clk),
    .D(_00660_),
    .RESET_B(net275),
    .Q(\u_rf.reg20_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12624_ (.CLK(clk),
    .D(_00661_),
    .RESET_B(net275),
    .Q(\u_rf.reg20_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12625_ (.CLK(clk),
    .D(_00662_),
    .RESET_B(net296),
    .Q(\u_rf.reg20_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12626_ (.CLK(clk),
    .D(_00663_),
    .RESET_B(net278),
    .Q(\u_rf.reg20_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12627_ (.CLK(clk),
    .D(_00664_),
    .RESET_B(net303),
    .Q(\u_rf.reg20_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12628_ (.CLK(clk),
    .D(_00665_),
    .RESET_B(net268),
    .Q(\u_rf.reg20_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12629_ (.CLK(clk),
    .D(_00666_),
    .RESET_B(net298),
    .Q(\u_rf.reg20_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12630_ (.CLK(clk),
    .D(_00667_),
    .RESET_B(net308),
    .Q(\u_rf.reg20_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12631_ (.CLK(clk),
    .D(_00668_),
    .RESET_B(net352),
    .Q(\u_rf.reg20_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12632_ (.CLK(clk),
    .D(_00669_),
    .RESET_B(net351),
    .Q(\u_rf.reg20_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12633_ (.CLK(clk),
    .D(_00670_),
    .RESET_B(net342),
    .Q(\u_rf.reg20_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12634_ (.CLK(clk),
    .D(_00671_),
    .RESET_B(net339),
    .Q(\u_rf.reg20_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12635_ (.CLK(clk),
    .D(_00672_),
    .RESET_B(net242),
    .Q(\u_rf.reg21_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12636_ (.CLK(clk),
    .D(_00673_),
    .RESET_B(net237),
    .Q(\u_rf.reg21_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12637_ (.CLK(clk),
    .D(_00674_),
    .RESET_B(net250),
    .Q(\u_rf.reg21_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12638_ (.CLK(clk),
    .D(_00675_),
    .RESET_B(net232),
    .Q(\u_rf.reg21_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12639_ (.CLK(clk),
    .D(_00676_),
    .RESET_B(net228),
    .Q(\u_rf.reg21_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12640_ (.CLK(clk),
    .D(_00677_),
    .RESET_B(net248),
    .Q(\u_rf.reg21_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12641_ (.CLK(clk),
    .D(_00678_),
    .RESET_B(net327),
    .Q(\u_rf.reg21_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12642_ (.CLK(clk),
    .D(_00679_),
    .RESET_B(net235),
    .Q(\u_rf.reg21_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12643_ (.CLK(clk),
    .D(_00680_),
    .RESET_B(net315),
    .Q(\u_rf.reg21_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12644_ (.CLK(clk),
    .D(_00681_),
    .RESET_B(net321),
    .Q(\u_rf.reg21_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12645_ (.CLK(clk),
    .D(_00682_),
    .RESET_B(net324),
    .Q(\u_rf.reg21_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12646_ (.CLK(clk),
    .D(_00683_),
    .RESET_B(net211),
    .Q(\u_rf.reg21_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12647_ (.CLK(clk),
    .D(_00684_),
    .RESET_B(net211),
    .Q(\u_rf.reg21_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12648_ (.CLK(clk),
    .D(_00685_),
    .RESET_B(net289),
    .Q(\u_rf.reg21_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12649_ (.CLK(clk),
    .D(_00686_),
    .RESET_B(net266),
    .Q(\u_rf.reg21_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12650_ (.CLK(clk),
    .D(_00687_),
    .RESET_B(net260),
    .Q(\u_rf.reg21_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12651_ (.CLK(clk),
    .D(_00688_),
    .RESET_B(net223),
    .Q(\u_rf.reg21_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12652_ (.CLK(clk),
    .D(_00689_),
    .RESET_B(net265),
    .Q(\u_rf.reg21_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12653_ (.CLK(clk),
    .D(_00690_),
    .RESET_B(net215),
    .Q(\u_rf.reg21_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12654_ (.CLK(clk),
    .D(_00691_),
    .RESET_B(net219),
    .Q(\u_rf.reg21_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12655_ (.CLK(clk),
    .D(_00692_),
    .RESET_B(net272),
    .Q(\u_rf.reg21_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12656_ (.CLK(clk),
    .D(_00693_),
    .RESET_B(net271),
    .Q(\u_rf.reg21_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12657_ (.CLK(clk),
    .D(_00694_),
    .RESET_B(net287),
    .Q(\u_rf.reg21_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12658_ (.CLK(clk),
    .D(_00695_),
    .RESET_B(net279),
    .Q(\u_rf.reg21_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12659_ (.CLK(clk),
    .D(_00696_),
    .RESET_B(net351),
    .Q(\u_rf.reg21_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12660_ (.CLK(clk),
    .D(_00697_),
    .RESET_B(net262),
    .Q(\u_rf.reg21_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12661_ (.CLK(clk),
    .D(_00698_),
    .RESET_B(net301),
    .Q(\u_rf.reg21_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12662_ (.CLK(clk),
    .D(_00699_),
    .RESET_B(net308),
    .Q(\u_rf.reg21_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12663_ (.CLK(clk),
    .D(_00700_),
    .RESET_B(net353),
    .Q(\u_rf.reg21_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12664_ (.CLK(clk),
    .D(_00701_),
    .RESET_B(net342),
    .Q(\u_rf.reg21_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12665_ (.CLK(clk),
    .D(_00702_),
    .RESET_B(net341),
    .Q(\u_rf.reg21_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12666_ (.CLK(clk),
    .D(_00703_),
    .RESET_B(net340),
    .Q(\u_rf.reg21_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12667_ (.CLK(clk),
    .D(_00704_),
    .RESET_B(net222),
    .Q(\u_rf.reg22_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12668_ (.CLK(clk),
    .D(_00705_),
    .RESET_B(net235),
    .Q(\u_rf.reg22_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12669_ (.CLK(clk),
    .D(_00706_),
    .RESET_B(net246),
    .Q(\u_rf.reg22_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12670_ (.CLK(clk),
    .D(_00707_),
    .RESET_B(net243),
    .Q(\u_rf.reg22_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12671_ (.CLK(clk),
    .D(_00708_),
    .RESET_B(net205),
    .Q(\u_rf.reg22_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12672_ (.CLK(clk),
    .D(_00709_),
    .RESET_B(net249),
    .Q(\u_rf.reg22_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12673_ (.CLK(clk),
    .D(_00710_),
    .RESET_B(net251),
    .Q(\u_rf.reg22_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12674_ (.CLK(clk),
    .D(_00711_),
    .RESET_B(net230),
    .Q(\u_rf.reg22_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12675_ (.CLK(clk),
    .D(_00712_),
    .RESET_B(net320),
    .Q(\u_rf.reg22_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12676_ (.CLK(clk),
    .D(_00713_),
    .RESET_B(net321),
    .Q(\u_rf.reg22_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12677_ (.CLK(clk),
    .D(_00714_),
    .RESET_B(net239),
    .Q(\u_rf.reg22_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12678_ (.CLK(clk),
    .D(_00715_),
    .RESET_B(net204),
    .Q(\u_rf.reg22_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12679_ (.CLK(clk),
    .D(_00716_),
    .RESET_B(net213),
    .Q(\u_rf.reg22_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12680_ (.CLK(clk),
    .D(_00717_),
    .RESET_B(net282),
    .Q(\u_rf.reg22_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12681_ (.CLK(clk),
    .D(_00718_),
    .RESET_B(net267),
    .Q(\u_rf.reg22_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12682_ (.CLK(clk),
    .D(_00719_),
    .RESET_B(net259),
    .Q(\u_rf.reg22_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12683_ (.CLK(clk),
    .D(_00720_),
    .RESET_B(net209),
    .Q(\u_rf.reg22_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12684_ (.CLK(clk),
    .D(_00721_),
    .RESET_B(net265),
    .Q(\u_rf.reg22_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12685_ (.CLK(clk),
    .D(_00722_),
    .RESET_B(net218),
    .Q(\u_rf.reg22_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12686_ (.CLK(clk),
    .D(_00723_),
    .RESET_B(net258),
    .Q(\u_rf.reg22_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12687_ (.CLK(clk),
    .D(_00724_),
    .RESET_B(net275),
    .Q(\u_rf.reg22_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12688_ (.CLK(clk),
    .D(_00725_),
    .RESET_B(net271),
    .Q(\u_rf.reg22_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12689_ (.CLK(clk),
    .D(_00726_),
    .RESET_B(net296),
    .Q(\u_rf.reg22_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12690_ (.CLK(clk),
    .D(_00727_),
    .RESET_B(net278),
    .Q(\u_rf.reg22_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12691_ (.CLK(clk),
    .D(_00728_),
    .RESET_B(net305),
    .Q(\u_rf.reg22_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12692_ (.CLK(clk),
    .D(_00729_),
    .RESET_B(net263),
    .Q(\u_rf.reg22_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12693_ (.CLK(clk),
    .D(_00730_),
    .RESET_B(net301),
    .Q(\u_rf.reg22_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12694_ (.CLK(clk),
    .D(_00731_),
    .RESET_B(net307),
    .Q(\u_rf.reg22_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12695_ (.CLK(clk),
    .D(_00732_),
    .RESET_B(net352),
    .Q(\u_rf.reg22_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12696_ (.CLK(clk),
    .D(_00733_),
    .RESET_B(net343),
    .Q(\u_rf.reg22_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12697_ (.CLK(clk),
    .D(_00734_),
    .RESET_B(net293),
    .Q(\u_rf.reg22_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12698_ (.CLK(clk),
    .D(_00735_),
    .RESET_B(net339),
    .Q(\u_rf.reg22_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12699_ (.CLK(clk),
    .D(_00736_),
    .RESET_B(net243),
    .Q(\u_rf.reg23_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12700_ (.CLK(clk),
    .D(_00737_),
    .RESET_B(net234),
    .Q(\u_rf.reg23_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12701_ (.CLK(clk),
    .D(_00738_),
    .RESET_B(net246),
    .Q(\u_rf.reg23_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12702_ (.CLK(clk),
    .D(_00739_),
    .RESET_B(net232),
    .Q(\u_rf.reg23_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12703_ (.CLK(clk),
    .D(_00740_),
    .RESET_B(net228),
    .Q(\u_rf.reg23_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12704_ (.CLK(clk),
    .D(_00741_),
    .RESET_B(net327),
    .Q(\u_rf.reg23_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12705_ (.CLK(clk),
    .D(_00742_),
    .RESET_B(net326),
    .Q(\u_rf.reg23_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12706_ (.CLK(clk),
    .D(_00743_),
    .RESET_B(net229),
    .Q(\u_rf.reg23_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12707_ (.CLK(clk),
    .D(_00744_),
    .RESET_B(net319),
    .Q(\u_rf.reg23_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12708_ (.CLK(clk),
    .D(_00745_),
    .RESET_B(net315),
    .Q(\u_rf.reg23_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12709_ (.CLK(clk),
    .D(_00746_),
    .RESET_B(net240),
    .Q(\u_rf.reg23_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12710_ (.CLK(clk),
    .D(_00747_),
    .RESET_B(net203),
    .Q(\u_rf.reg23_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12711_ (.CLK(clk),
    .D(_00748_),
    .RESET_B(net214),
    .Q(\u_rf.reg23_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12712_ (.CLK(clk),
    .D(_00749_),
    .RESET_B(net291),
    .Q(\u_rf.reg23_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12713_ (.CLK(clk),
    .D(_00750_),
    .RESET_B(net284),
    .Q(\u_rf.reg23_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12714_ (.CLK(clk),
    .D(_00751_),
    .RESET_B(net262),
    .Q(\u_rf.reg23_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12715_ (.CLK(clk),
    .D(_00752_),
    .RESET_B(net207),
    .Q(\u_rf.reg23_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12716_ (.CLK(clk),
    .D(_00753_),
    .RESET_B(net224),
    .Q(\u_rf.reg23_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12717_ (.CLK(clk),
    .D(_00754_),
    .RESET_B(net217),
    .Q(\u_rf.reg23_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12718_ (.CLK(clk),
    .D(_00755_),
    .RESET_B(net218),
    .Q(\u_rf.reg23_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12719_ (.CLK(clk),
    .D(_00756_),
    .RESET_B(net275),
    .Q(\u_rf.reg23_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12720_ (.CLK(clk),
    .D(_00757_),
    .RESET_B(net268),
    .Q(\u_rf.reg23_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12721_ (.CLK(clk),
    .D(_00758_),
    .RESET_B(net293),
    .Q(\u_rf.reg23_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12722_ (.CLK(clk),
    .D(_00759_),
    .RESET_B(net279),
    .Q(\u_rf.reg23_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12723_ (.CLK(clk),
    .D(_00760_),
    .RESET_B(net351),
    .Q(\u_rf.reg23_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12724_ (.CLK(clk),
    .D(_00761_),
    .RESET_B(net267),
    .Q(\u_rf.reg23_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12725_ (.CLK(clk),
    .D(_00762_),
    .RESET_B(net295),
    .Q(\u_rf.reg23_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12726_ (.CLK(clk),
    .D(_00763_),
    .RESET_B(net309),
    .Q(\u_rf.reg23_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12727_ (.CLK(clk),
    .D(_00764_),
    .RESET_B(net352),
    .Q(\u_rf.reg23_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12728_ (.CLK(clk),
    .D(_00765_),
    .RESET_B(net351),
    .Q(\u_rf.reg23_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12729_ (.CLK(clk),
    .D(_00766_),
    .RESET_B(net342),
    .Q(\u_rf.reg23_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12730_ (.CLK(clk),
    .D(_00767_),
    .RESET_B(net341),
    .Q(\u_rf.reg23_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12731_ (.CLK(clk),
    .D(_00768_),
    .RESET_B(net222),
    .Q(\u_rf.reg24_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12732_ (.CLK(clk),
    .D(_00769_),
    .RESET_B(net237),
    .Q(\u_rf.reg24_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12733_ (.CLK(clk),
    .D(_00770_),
    .RESET_B(net281),
    .Q(\u_rf.reg24_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12734_ (.CLK(clk),
    .D(_00771_),
    .RESET_B(net209),
    .Q(\u_rf.reg24_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12735_ (.CLK(clk),
    .D(_00772_),
    .RESET_B(net206),
    .Q(\u_rf.reg24_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12736_ (.CLK(clk),
    .D(_00773_),
    .RESET_B(net327),
    .Q(\u_rf.reg24_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12737_ (.CLK(clk),
    .D(_00774_),
    .RESET_B(net325),
    .Q(\u_rf.reg24_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12738_ (.CLK(clk),
    .D(_00775_),
    .RESET_B(net230),
    .Q(\u_rf.reg24_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12739_ (.CLK(clk),
    .D(_00776_),
    .RESET_B(net320),
    .Q(\u_rf.reg24_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12740_ (.CLK(clk),
    .D(_00777_),
    .RESET_B(net317),
    .Q(\u_rf.reg24_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12741_ (.CLK(clk),
    .D(_00778_),
    .RESET_B(net247),
    .Q(\u_rf.reg24_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12742_ (.CLK(clk),
    .D(_00779_),
    .RESET_B(net203),
    .Q(\u_rf.reg24_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12743_ (.CLK(clk),
    .D(_00780_),
    .RESET_B(net212),
    .Q(\u_rf.reg24_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12744_ (.CLK(clk),
    .D(_00781_),
    .RESET_B(net290),
    .Q(\u_rf.reg24_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12745_ (.CLK(clk),
    .D(_00782_),
    .RESET_B(net286),
    .Q(\u_rf.reg24_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12746_ (.CLK(clk),
    .D(_00783_),
    .RESET_B(net261),
    .Q(\u_rf.reg24_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12747_ (.CLK(clk),
    .D(_00784_),
    .RESET_B(net208),
    .Q(\u_rf.reg24_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12748_ (.CLK(clk),
    .D(_00785_),
    .RESET_B(net265),
    .Q(\u_rf.reg24_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12749_ (.CLK(clk),
    .D(_00786_),
    .RESET_B(net216),
    .Q(\u_rf.reg24_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12750_ (.CLK(clk),
    .D(_00787_),
    .RESET_B(net256),
    .Q(\u_rf.reg24_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12751_ (.CLK(clk),
    .D(_00788_),
    .RESET_B(net272),
    .Q(\u_rf.reg24_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12752_ (.CLK(clk),
    .D(_00789_),
    .RESET_B(net271),
    .Q(\u_rf.reg24_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12753_ (.CLK(clk),
    .D(_00790_),
    .RESET_B(net286),
    .Q(\u_rf.reg24_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12754_ (.CLK(clk),
    .D(_00791_),
    .RESET_B(net277),
    .Q(\u_rf.reg24_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12755_ (.CLK(clk),
    .D(_00792_),
    .RESET_B(net304),
    .Q(\u_rf.reg24_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12756_ (.CLK(clk),
    .D(_00793_),
    .RESET_B(net262),
    .Q(\u_rf.reg24_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12757_ (.CLK(clk),
    .D(_00794_),
    .RESET_B(net300),
    .Q(\u_rf.reg24_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12758_ (.CLK(clk),
    .D(_00795_),
    .RESET_B(net307),
    .Q(\u_rf.reg24_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12759_ (.CLK(clk),
    .D(_00796_),
    .RESET_B(net352),
    .Q(\u_rf.reg24_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12760_ (.CLK(clk),
    .D(_00797_),
    .RESET_B(net343),
    .Q(\u_rf.reg24_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12761_ (.CLK(clk),
    .D(_00798_),
    .RESET_B(net292),
    .Q(\u_rf.reg24_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12762_ (.CLK(clk),
    .D(_00799_),
    .RESET_B(net290),
    .Q(\u_rf.reg24_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12763_ (.CLK(clk),
    .D(_00800_),
    .RESET_B(net244),
    .Q(\u_rf.reg25_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12764_ (.CLK(clk),
    .D(_00801_),
    .RESET_B(net238),
    .Q(\u_rf.reg25_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12765_ (.CLK(clk),
    .D(_00802_),
    .RESET_B(net281),
    .Q(\u_rf.reg25_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12766_ (.CLK(clk),
    .D(_00803_),
    .RESET_B(net232),
    .Q(\u_rf.reg25_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12767_ (.CLK(clk),
    .D(_00804_),
    .RESET_B(net228),
    .Q(\u_rf.reg25_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12768_ (.CLK(clk),
    .D(_00805_),
    .RESET_B(net249),
    .Q(\u_rf.reg25_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12769_ (.CLK(clk),
    .D(_00806_),
    .RESET_B(net251),
    .Q(\u_rf.reg25_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12770_ (.CLK(clk),
    .D(_00807_),
    .RESET_B(net235),
    .Q(\u_rf.reg25_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12771_ (.CLK(clk),
    .D(_00808_),
    .RESET_B(net313),
    .Q(\u_rf.reg25_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12772_ (.CLK(clk),
    .D(_00809_),
    .RESET_B(net316),
    .Q(\u_rf.reg25_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12773_ (.CLK(clk),
    .D(_00810_),
    .RESET_B(net247),
    .Q(\u_rf.reg25_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12774_ (.CLK(clk),
    .D(_00811_),
    .RESET_B(net204),
    .Q(\u_rf.reg25_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12775_ (.CLK(clk),
    .D(_00812_),
    .RESET_B(net211),
    .Q(\u_rf.reg25_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12776_ (.CLK(clk),
    .D(_00813_),
    .RESET_B(net289),
    .Q(\u_rf.reg25_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12777_ (.CLK(clk),
    .D(_00814_),
    .RESET_B(net283),
    .Q(\u_rf.reg25_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12778_ (.CLK(clk),
    .D(_00815_),
    .RESET_B(net260),
    .Q(\u_rf.reg25_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12779_ (.CLK(clk),
    .D(_00816_),
    .RESET_B(net223),
    .Q(\u_rf.reg25_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12780_ (.CLK(clk),
    .D(_00817_),
    .RESET_B(net280),
    .Q(\u_rf.reg25_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12781_ (.CLK(clk),
    .D(_00818_),
    .RESET_B(net217),
    .Q(\u_rf.reg25_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12782_ (.CLK(clk),
    .D(_00819_),
    .RESET_B(net257),
    .Q(\u_rf.reg25_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12783_ (.CLK(clk),
    .D(_00820_),
    .RESET_B(net272),
    .Q(\u_rf.reg25_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12784_ (.CLK(clk),
    .D(_00821_),
    .RESET_B(net271),
    .Q(\u_rf.reg25_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12785_ (.CLK(clk),
    .D(_00822_),
    .RESET_B(net287),
    .Q(\u_rf.reg25_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12786_ (.CLK(clk),
    .D(_00823_),
    .RESET_B(net274),
    .Q(\u_rf.reg25_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12787_ (.CLK(clk),
    .D(_00824_),
    .RESET_B(net350),
    .Q(\u_rf.reg25_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12788_ (.CLK(clk),
    .D(_00825_),
    .RESET_B(net263),
    .Q(\u_rf.reg25_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12789_ (.CLK(clk),
    .D(_00826_),
    .RESET_B(net301),
    .Q(\u_rf.reg25_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12790_ (.CLK(clk),
    .D(_00827_),
    .RESET_B(net306),
    .Q(\u_rf.reg25_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12791_ (.CLK(clk),
    .D(_00828_),
    .RESET_B(net353),
    .Q(\u_rf.reg25_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12792_ (.CLK(clk),
    .D(_00829_),
    .RESET_B(net349),
    .Q(\u_rf.reg25_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12793_ (.CLK(clk),
    .D(_00830_),
    .RESET_B(net346),
    .Q(\u_rf.reg25_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12794_ (.CLK(clk),
    .D(_00831_),
    .RESET_B(net340),
    .Q(\u_rf.reg25_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12795_ (.CLK(clk),
    .D(_00832_),
    .RESET_B(net248),
    .Q(\u_rf.reg26_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12796_ (.CLK(clk),
    .D(_00833_),
    .RESET_B(net240),
    .Q(\u_rf.reg26_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12797_ (.CLK(clk),
    .D(_00834_),
    .RESET_B(net250),
    .Q(\u_rf.reg26_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12798_ (.CLK(clk),
    .D(_00835_),
    .RESET_B(net241),
    .Q(\u_rf.reg26_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12799_ (.CLK(clk),
    .D(_00836_),
    .RESET_B(net228),
    .Q(\u_rf.reg26_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12800_ (.CLK(clk),
    .D(_00837_),
    .RESET_B(net330),
    .Q(\u_rf.reg26_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12801_ (.CLK(clk),
    .D(_00838_),
    .RESET_B(net325),
    .Q(\u_rf.reg26_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12802_ (.CLK(clk),
    .D(_00839_),
    .RESET_B(net235),
    .Q(\u_rf.reg26_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12803_ (.CLK(clk),
    .D(_00840_),
    .RESET_B(net320),
    .Q(\u_rf.reg26_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12804_ (.CLK(clk),
    .D(_00841_),
    .RESET_B(net322),
    .Q(\u_rf.reg26_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12805_ (.CLK(clk),
    .D(_00842_),
    .RESET_B(net324),
    .Q(\u_rf.reg26_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12806_ (.CLK(clk),
    .D(_00843_),
    .RESET_B(net213),
    .Q(\u_rf.reg26_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12807_ (.CLK(clk),
    .D(_00844_),
    .RESET_B(net213),
    .Q(\u_rf.reg26_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12808_ (.CLK(clk),
    .D(_00845_),
    .RESET_B(net290),
    .Q(\u_rf.reg26_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12809_ (.CLK(clk),
    .D(_00846_),
    .RESET_B(net283),
    .Q(\u_rf.reg26_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12810_ (.CLK(clk),
    .D(_00847_),
    .RESET_B(net259),
    .Q(\u_rf.reg26_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12811_ (.CLK(clk),
    .D(_00848_),
    .RESET_B(net222),
    .Q(\u_rf.reg26_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12812_ (.CLK(clk),
    .D(_00849_),
    .RESET_B(net280),
    .Q(\u_rf.reg26_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12813_ (.CLK(clk),
    .D(_00850_),
    .RESET_B(net217),
    .Q(\u_rf.reg26_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12814_ (.CLK(clk),
    .D(_00851_),
    .RESET_B(net218),
    .Q(\u_rf.reg26_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12815_ (.CLK(clk),
    .D(_00852_),
    .RESET_B(net276),
    .Q(\u_rf.reg26_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12816_ (.CLK(clk),
    .D(_00853_),
    .RESET_B(net275),
    .Q(\u_rf.reg26_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12817_ (.CLK(clk),
    .D(_00854_),
    .RESET_B(net293),
    .Q(\u_rf.reg26_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12818_ (.CLK(clk),
    .D(_00855_),
    .RESET_B(net278),
    .Q(\u_rf.reg26_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12819_ (.CLK(clk),
    .D(_00856_),
    .RESET_B(net356),
    .Q(\u_rf.reg26_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12820_ (.CLK(clk),
    .D(_00857_),
    .RESET_B(net285),
    .Q(\u_rf.reg26_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12821_ (.CLK(clk),
    .D(_00858_),
    .RESET_B(net297),
    .Q(\u_rf.reg26_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12822_ (.CLK(clk),
    .D(_00859_),
    .RESET_B(net358),
    .Q(\u_rf.reg26_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12823_ (.CLK(clk),
    .D(_00860_),
    .RESET_B(net359),
    .Q(\u_rf.reg26_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12824_ (.CLK(clk),
    .D(_00861_),
    .RESET_B(net355),
    .Q(\u_rf.reg26_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12825_ (.CLK(clk),
    .D(_00862_),
    .RESET_B(net346),
    .Q(\u_rf.reg26_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12826_ (.CLK(clk),
    .D(_00863_),
    .RESET_B(net344),
    .Q(\u_rf.reg26_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12827_ (.CLK(clk),
    .D(_00864_),
    .RESET_B(net224),
    .Q(\u_rf.reg27_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12828_ (.CLK(clk),
    .D(_00865_),
    .RESET_B(net237),
    .Q(\u_rf.reg27_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12829_ (.CLK(clk),
    .D(_00866_),
    .RESET_B(net244),
    .Q(\u_rf.reg27_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12830_ (.CLK(clk),
    .D(_00867_),
    .RESET_B(net228),
    .Q(\u_rf.reg27_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12831_ (.CLK(clk),
    .D(_00868_),
    .RESET_B(net206),
    .Q(\u_rf.reg27_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12832_ (.CLK(clk),
    .D(_00869_),
    .RESET_B(net249),
    .Q(\u_rf.reg27_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12833_ (.CLK(clk),
    .D(_00870_),
    .RESET_B(net326),
    .Q(\u_rf.reg27_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12834_ (.CLK(clk),
    .D(_00871_),
    .RESET_B(net230),
    .Q(\u_rf.reg27_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12835_ (.CLK(clk),
    .D(_00872_),
    .RESET_B(net312),
    .Q(\u_rf.reg27_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12836_ (.CLK(clk),
    .D(_00873_),
    .RESET_B(net316),
    .Q(\u_rf.reg27_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12837_ (.CLK(clk),
    .D(_00874_),
    .RESET_B(net231),
    .Q(\u_rf.reg27_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12838_ (.CLK(clk),
    .D(_00875_),
    .RESET_B(net204),
    .Q(\u_rf.reg27_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12839_ (.CLK(clk),
    .D(_00876_),
    .RESET_B(net214),
    .Q(\u_rf.reg27_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12840_ (.CLK(clk),
    .D(_00877_),
    .RESET_B(net286),
    .Q(\u_rf.reg27_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12841_ (.CLK(clk),
    .D(_00878_),
    .RESET_B(net284),
    .Q(\u_rf.reg27_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12842_ (.CLK(clk),
    .D(_00879_),
    .RESET_B(net259),
    .Q(\u_rf.reg27_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12843_ (.CLK(clk),
    .D(_00880_),
    .RESET_B(net207),
    .Q(\u_rf.reg27_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12844_ (.CLK(clk),
    .D(_00881_),
    .RESET_B(net225),
    .Q(\u_rf.reg27_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12845_ (.CLK(clk),
    .D(_00882_),
    .RESET_B(net224),
    .Q(\u_rf.reg27_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12846_ (.CLK(clk),
    .D(_00883_),
    .RESET_B(net218),
    .Q(\u_rf.reg27_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12847_ (.CLK(clk),
    .D(_00884_),
    .RESET_B(net273),
    .Q(\u_rf.reg27_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12848_ (.CLK(clk),
    .D(_00885_),
    .RESET_B(net264),
    .Q(\u_rf.reg27_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12849_ (.CLK(clk),
    .D(_00886_),
    .RESET_B(net294),
    .Q(\u_rf.reg27_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12850_ (.CLK(clk),
    .D(_00887_),
    .RESET_B(net279),
    .Q(\u_rf.reg27_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12851_ (.CLK(clk),
    .D(_00888_),
    .RESET_B(net351),
    .Q(\u_rf.reg27_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12852_ (.CLK(clk),
    .D(_00889_),
    .RESET_B(net264),
    .Q(\u_rf.reg27_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12853_ (.CLK(clk),
    .D(_00890_),
    .RESET_B(net299),
    .Q(\u_rf.reg27_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12854_ (.CLK(clk),
    .D(_00891_),
    .RESET_B(net306),
    .Q(\u_rf.reg27_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12855_ (.CLK(clk),
    .D(_00892_),
    .RESET_B(net354),
    .Q(\u_rf.reg27_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12856_ (.CLK(clk),
    .D(_00893_),
    .RESET_B(net304),
    .Q(\u_rf.reg27_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12857_ (.CLK(clk),
    .D(_00894_),
    .RESET_B(net341),
    .Q(\u_rf.reg27_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12858_ (.CLK(clk),
    .D(_00895_),
    .RESET_B(net341),
    .Q(\u_rf.reg27_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12859_ (.CLK(clk),
    .D(_00896_),
    .RESET_B(net242),
    .Q(\u_rf.reg28_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12860_ (.CLK(clk),
    .D(_00897_),
    .RESET_B(net316),
    .Q(\u_rf.reg28_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12861_ (.CLK(clk),
    .D(_00898_),
    .RESET_B(net250),
    .Q(\u_rf.reg28_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12862_ (.CLK(clk),
    .D(_00899_),
    .RESET_B(net241),
    .Q(\u_rf.reg28_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12863_ (.CLK(clk),
    .D(_00900_),
    .RESET_B(net231),
    .Q(\u_rf.reg28_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12864_ (.CLK(clk),
    .D(_00901_),
    .RESET_B(net327),
    .Q(\u_rf.reg28_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12865_ (.CLK(clk),
    .D(_00902_),
    .RESET_B(net325),
    .Q(\u_rf.reg28_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12866_ (.CLK(clk),
    .D(_00903_),
    .RESET_B(net239),
    .Q(\u_rf.reg28_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12867_ (.CLK(clk),
    .D(_00904_),
    .RESET_B(net321),
    .Q(\u_rf.reg28_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12868_ (.CLK(clk),
    .D(_00905_),
    .RESET_B(net317),
    .Q(\u_rf.reg28_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12869_ (.CLK(clk),
    .D(_00906_),
    .RESET_B(net249),
    .Q(\u_rf.reg28_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12870_ (.CLK(clk),
    .D(_00907_),
    .RESET_B(net213),
    .Q(\u_rf.reg28_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12871_ (.CLK(clk),
    .D(_00908_),
    .RESET_B(net223),
    .Q(\u_rf.reg28_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12872_ (.CLK(clk),
    .D(_00909_),
    .RESET_B(net288),
    .Q(\u_rf.reg28_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12873_ (.CLK(clk),
    .D(_00910_),
    .RESET_B(net283),
    .Q(\u_rf.reg28_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12874_ (.CLK(clk),
    .D(_00911_),
    .RESET_B(net266),
    .Q(\u_rf.reg28_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12875_ (.CLK(clk),
    .D(_00912_),
    .RESET_B(net223),
    .Q(\u_rf.reg28_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12876_ (.CLK(clk),
    .D(_00913_),
    .RESET_B(net281),
    .Q(\u_rf.reg28_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12877_ (.CLK(clk),
    .D(_00914_),
    .RESET_B(net224),
    .Q(\u_rf.reg28_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12878_ (.CLK(clk),
    .D(_00915_),
    .RESET_B(net226),
    .Q(\u_rf.reg28_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12879_ (.CLK(clk),
    .D(_00916_),
    .RESET_B(net295),
    .Q(\u_rf.reg28_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12880_ (.CLK(clk),
    .D(_00917_),
    .RESET_B(net294),
    .Q(\u_rf.reg28_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12881_ (.CLK(clk),
    .D(_00918_),
    .RESET_B(net302),
    .Q(\u_rf.reg28_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12882_ (.CLK(clk),
    .D(_00919_),
    .RESET_B(net298),
    .Q(\u_rf.reg28_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12883_ (.CLK(clk),
    .D(_00920_),
    .RESET_B(net356),
    .Q(\u_rf.reg28_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12884_ (.CLK(clk),
    .D(_00921_),
    .RESET_B(net285),
    .Q(\u_rf.reg28_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12885_ (.CLK(clk),
    .D(_00922_),
    .RESET_B(net303),
    .Q(\u_rf.reg28_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12886_ (.CLK(clk),
    .D(_00923_),
    .RESET_B(net359),
    .Q(\u_rf.reg28_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12887_ (.CLK(clk),
    .D(_00924_),
    .RESET_B(net359),
    .Q(\u_rf.reg28_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12888_ (.CLK(clk),
    .D(_00925_),
    .RESET_B(net355),
    .Q(\u_rf.reg28_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12889_ (.CLK(clk),
    .D(_00926_),
    .RESET_B(net346),
    .Q(\u_rf.reg28_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12890_ (.CLK(clk),
    .D(_00927_),
    .RESET_B(net344),
    .Q(\u_rf.reg28_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12891_ (.CLK(clk),
    .D(_00928_),
    .RESET_B(net221),
    .Q(\u_rf.reg29_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12892_ (.CLK(clk),
    .D(_00929_),
    .RESET_B(net236),
    .Q(\u_rf.reg29_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12893_ (.CLK(clk),
    .D(_00930_),
    .RESET_B(net250),
    .Q(\u_rf.reg29_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12894_ (.CLK(clk),
    .D(_00931_),
    .RESET_B(net221),
    .Q(\u_rf.reg29_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12895_ (.CLK(clk),
    .D(_00932_),
    .RESET_B(net227),
    .Q(\u_rf.reg29_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12896_ (.CLK(clk),
    .D(_00933_),
    .RESET_B(net324),
    .Q(\u_rf.reg29_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12897_ (.CLK(clk),
    .D(_00934_),
    .RESET_B(net252),
    .Q(\u_rf.reg29_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12898_ (.CLK(clk),
    .D(_00935_),
    .RESET_B(net229),
    .Q(\u_rf.reg29_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12899_ (.CLK(clk),
    .D(_00936_),
    .RESET_B(net314),
    .Q(\u_rf.reg29_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12900_ (.CLK(clk),
    .D(_00937_),
    .RESET_B(net315),
    .Q(\u_rf.reg29_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12901_ (.CLK(clk),
    .D(_00938_),
    .RESET_B(net240),
    .Q(\u_rf.reg29_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12902_ (.CLK(clk),
    .D(_00939_),
    .RESET_B(net204),
    .Q(\u_rf.reg29_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12903_ (.CLK(clk),
    .D(_00940_),
    .RESET_B(net213),
    .Q(\u_rf.reg29_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12904_ (.CLK(clk),
    .D(_00941_),
    .RESET_B(net286),
    .Q(\u_rf.reg29_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12905_ (.CLK(clk),
    .D(_00942_),
    .RESET_B(net267),
    .Q(\u_rf.reg29_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12906_ (.CLK(clk),
    .D(_00943_),
    .RESET_B(net259),
    .Q(\u_rf.reg29_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12907_ (.CLK(clk),
    .D(_00944_),
    .RESET_B(net209),
    .Q(\u_rf.reg29_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12908_ (.CLK(clk),
    .D(_00945_),
    .RESET_B(net225),
    .Q(\u_rf.reg29_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12909_ (.CLK(clk),
    .D(_00946_),
    .RESET_B(net226),
    .Q(\u_rf.reg29_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12910_ (.CLK(clk),
    .D(_00947_),
    .RESET_B(net258),
    .Q(\u_rf.reg29_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12911_ (.CLK(clk),
    .D(_00948_),
    .RESET_B(net272),
    .Q(\u_rf.reg29_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12912_ (.CLK(clk),
    .D(_00949_),
    .RESET_B(net271),
    .Q(\u_rf.reg29_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12913_ (.CLK(clk),
    .D(_00950_),
    .RESET_B(net285),
    .Q(\u_rf.reg29_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12914_ (.CLK(clk),
    .D(_00951_),
    .RESET_B(net279),
    .Q(\u_rf.reg29_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12915_ (.CLK(clk),
    .D(_00952_),
    .RESET_B(net351),
    .Q(\u_rf.reg29_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12916_ (.CLK(clk),
    .D(_00953_),
    .RESET_B(net268),
    .Q(\u_rf.reg29_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12917_ (.CLK(clk),
    .D(_00954_),
    .RESET_B(net301),
    .Q(\u_rf.reg29_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12918_ (.CLK(clk),
    .D(_00955_),
    .RESET_B(net309),
    .Q(\u_rf.reg29_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12919_ (.CLK(clk),
    .D(_00956_),
    .RESET_B(net354),
    .Q(\u_rf.reg29_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12920_ (.CLK(clk),
    .D(_00957_),
    .RESET_B(net349),
    .Q(\u_rf.reg29_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12921_ (.CLK(clk),
    .D(_00958_),
    .RESET_B(net342),
    .Q(\u_rf.reg29_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12922_ (.CLK(clk),
    .D(_00959_),
    .RESET_B(net339),
    .Q(\u_rf.reg29_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12923_ (.CLK(clk),
    .D(_00960_),
    .RESET_B(net242),
    .Q(\u_rf.reg30_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12924_ (.CLK(clk),
    .D(_00961_),
    .RESET_B(net240),
    .Q(\u_rf.reg30_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12925_ (.CLK(clk),
    .D(_00962_),
    .RESET_B(net252),
    .Q(\u_rf.reg30_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12926_ (.CLK(clk),
    .D(_00963_),
    .RESET_B(net231),
    .Q(\u_rf.reg30_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12927_ (.CLK(clk),
    .D(_00964_),
    .RESET_B(net233),
    .Q(\u_rf.reg30_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12928_ (.CLK(clk),
    .D(_00965_),
    .RESET_B(net323),
    .Q(\u_rf.reg30_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12929_ (.CLK(clk),
    .D(_00966_),
    .RESET_B(net327),
    .Q(\u_rf.reg30_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12930_ (.CLK(clk),
    .D(_00967_),
    .RESET_B(net234),
    .Q(\u_rf.reg30_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12931_ (.CLK(clk),
    .D(_00968_),
    .RESET_B(net319),
    .Q(\u_rf.reg30_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12932_ (.CLK(clk),
    .D(_00969_),
    .RESET_B(net320),
    .Q(\u_rf.reg30_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12933_ (.CLK(clk),
    .D(_00970_),
    .RESET_B(net249),
    .Q(\u_rf.reg30_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12934_ (.CLK(clk),
    .D(_00971_),
    .RESET_B(net210),
    .Q(\u_rf.reg30_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12935_ (.CLK(clk),
    .D(_00972_),
    .RESET_B(net214),
    .Q(\u_rf.reg30_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12936_ (.CLK(clk),
    .D(_00973_),
    .RESET_B(net291),
    .Q(\u_rf.reg30_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12937_ (.CLK(clk),
    .D(_00974_),
    .RESET_B(net284),
    .Q(\u_rf.reg30_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12938_ (.CLK(clk),
    .D(_00975_),
    .RESET_B(net262),
    .Q(\u_rf.reg30_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12939_ (.CLK(clk),
    .D(_00976_),
    .RESET_B(net205),
    .Q(\u_rf.reg30_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12940_ (.CLK(clk),
    .D(_00977_),
    .RESET_B(net224),
    .Q(\u_rf.reg30_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12941_ (.CLK(clk),
    .D(_00978_),
    .RESET_B(net226),
    .Q(\u_rf.reg30_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12942_ (.CLK(clk),
    .D(_00979_),
    .RESET_B(net218),
    .Q(\u_rf.reg30_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12943_ (.CLK(clk),
    .D(_00980_),
    .RESET_B(net295),
    .Q(\u_rf.reg30_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12944_ (.CLK(clk),
    .D(_00981_),
    .RESET_B(net285),
    .Q(\u_rf.reg30_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12945_ (.CLK(clk),
    .D(_00982_),
    .RESET_B(net296),
    .Q(\u_rf.reg30_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12946_ (.CLK(clk),
    .D(_00983_),
    .RESET_B(net299),
    .Q(\u_rf.reg30_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12947_ (.CLK(clk),
    .D(_00984_),
    .RESET_B(net303),
    .Q(\u_rf.reg30_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12948_ (.CLK(clk),
    .D(_00985_),
    .RESET_B(net284),
    .Q(\u_rf.reg30_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12949_ (.CLK(clk),
    .D(_00986_),
    .RESET_B(net297),
    .Q(\u_rf.reg30_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12950_ (.CLK(clk),
    .D(_00987_),
    .RESET_B(net309),
    .Q(\u_rf.reg30_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12951_ (.CLK(clk),
    .D(_00988_),
    .RESET_B(net354),
    .Q(\u_rf.reg30_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12952_ (.CLK(clk),
    .D(_00989_),
    .RESET_B(net349),
    .Q(\u_rf.reg30_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12953_ (.CLK(clk),
    .D(_00990_),
    .RESET_B(net341),
    .Q(\u_rf.reg30_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12954_ (.CLK(clk),
    .D(_00991_),
    .RESET_B(net340),
    .Q(\u_rf.reg30_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12955_ (.CLK(clk),
    .D(_00992_),
    .RESET_B(net242),
    .Q(\u_rf.reg31_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12956_ (.CLK(clk),
    .D(_00993_),
    .RESET_B(net238),
    .Q(\u_rf.reg31_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12957_ (.CLK(clk),
    .D(_00994_),
    .RESET_B(net246),
    .Q(\u_rf.reg31_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12958_ (.CLK(clk),
    .D(_00995_),
    .RESET_B(net232),
    .Q(\u_rf.reg31_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12959_ (.CLK(clk),
    .D(_00996_),
    .RESET_B(net230),
    .Q(\u_rf.reg31_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12960_ (.CLK(clk),
    .D(_00997_),
    .RESET_B(net324),
    .Q(\u_rf.reg31_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12961_ (.CLK(clk),
    .D(_00998_),
    .RESET_B(net326),
    .Q(\u_rf.reg31_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12962_ (.CLK(clk),
    .D(_00999_),
    .RESET_B(net235),
    .Q(\u_rf.reg31_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12963_ (.CLK(clk),
    .D(_01000_),
    .RESET_B(net315),
    .Q(\u_rf.reg31_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12964_ (.CLK(clk),
    .D(_01001_),
    .RESET_B(net315),
    .Q(\u_rf.reg31_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12965_ (.CLK(clk),
    .D(_01002_),
    .RESET_B(net240),
    .Q(\u_rf.reg31_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12966_ (.CLK(clk),
    .D(_01003_),
    .RESET_B(net203),
    .Q(\u_rf.reg31_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12967_ (.CLK(clk),
    .D(_01004_),
    .RESET_B(net214),
    .Q(\u_rf.reg31_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12968_ (.CLK(clk),
    .D(_01005_),
    .RESET_B(net289),
    .Q(\u_rf.reg31_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12969_ (.CLK(clk),
    .D(_01006_),
    .RESET_B(net282),
    .Q(\u_rf.reg31_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12970_ (.CLK(clk),
    .D(_01007_),
    .RESET_B(net259),
    .Q(\u_rf.reg31_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12971_ (.CLK(clk),
    .D(_01008_),
    .RESET_B(net205),
    .Q(\u_rf.reg31_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12972_ (.CLK(clk),
    .D(_01009_),
    .RESET_B(net246),
    .Q(\u_rf.reg31_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12973_ (.CLK(clk),
    .D(_01010_),
    .RESET_B(net224),
    .Q(\u_rf.reg31_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12974_ (.CLK(clk),
    .D(_01011_),
    .RESET_B(net258),
    .Q(\u_rf.reg31_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12975_ (.CLK(clk),
    .D(_01012_),
    .RESET_B(net294),
    .Q(\u_rf.reg31_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12976_ (.CLK(clk),
    .D(_01013_),
    .RESET_B(net294),
    .Q(\u_rf.reg31_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12977_ (.CLK(clk),
    .D(_01014_),
    .RESET_B(net294),
    .Q(\u_rf.reg31_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12978_ (.CLK(clk),
    .D(_01015_),
    .RESET_B(net299),
    .Q(\u_rf.reg31_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12979_ (.CLK(clk),
    .D(_01016_),
    .RESET_B(net303),
    .Q(\u_rf.reg31_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12980_ (.CLK(clk),
    .D(_01017_),
    .RESET_B(net285),
    .Q(\u_rf.reg31_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12981_ (.CLK(clk),
    .D(_01018_),
    .RESET_B(net298),
    .Q(\u_rf.reg31_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12982_ (.CLK(clk),
    .D(_01019_),
    .RESET_B(net309),
    .Q(\u_rf.reg31_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12983_ (.CLK(clk),
    .D(_01020_),
    .RESET_B(net352),
    .Q(\u_rf.reg31_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12984_ (.CLK(clk),
    .D(_01021_),
    .RESET_B(net351),
    .Q(\u_rf.reg31_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12985_ (.CLK(clk),
    .D(_01022_),
    .RESET_B(net346),
    .Q(\u_rf.reg31_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12986_ (.CLK(clk),
    .D(_01023_),
    .RESET_B(net340),
    .Q(\u_rf.reg31_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12987_ (.CLK(clk),
    .D(_01024_),
    .Q(\u_decod.branch_imm_q_o[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12988_ (.CLK(clk),
    .D(_01025_),
    .Q(\u_decod.branch_imm_q_o[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12989_ (.CLK(clk),
    .D(_01026_),
    .Q(\u_decod.branch_imm_q_o[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clk),
    .D(_01027_),
    .Q(\u_decod.branch_imm_q_o[3] ));
 sky130_fd_sc_hd__dfxtp_2 _12991_ (.CLK(clk),
    .D(_01028_),
    .Q(\u_decod.branch_imm_q_o[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clk),
    .D(_01029_),
    .Q(\u_decod.branch_imm_q_o[5] ));
 sky130_fd_sc_hd__dfxtp_2 _12993_ (.CLK(clk),
    .D(_01030_),
    .Q(\u_decod.branch_imm_q_o[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clk),
    .D(_01031_),
    .Q(\u_decod.branch_imm_q_o[7] ));
 sky130_fd_sc_hd__dfxtp_2 _12995_ (.CLK(clk),
    .D(_01032_),
    .Q(\u_decod.branch_imm_q_o[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clk),
    .D(_01033_),
    .Q(\u_decod.branch_imm_q_o[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12997_ (.CLK(clk),
    .D(_01034_),
    .Q(\u_decod.branch_imm_q_o[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12998_ (.CLK(clk),
    .D(_01035_),
    .Q(\u_decod.branch_imm_q_o[11] ));
 sky130_fd_sc_hd__dfxtp_2 _12999_ (.CLK(clk),
    .D(_01036_),
    .Q(\u_decod.branch_imm_q_o[12] ));
 sky130_fd_sc_hd__dfxtp_2 _13000_ (.CLK(clk),
    .D(_01037_),
    .Q(\u_decod.branch_imm_q_o[13] ));
 sky130_fd_sc_hd__dfxtp_2 _13001_ (.CLK(clk),
    .D(_01038_),
    .Q(\u_decod.branch_imm_q_o[14] ));
 sky130_fd_sc_hd__dfxtp_2 _13002_ (.CLK(clk),
    .D(_01039_),
    .Q(\u_decod.branch_imm_q_o[15] ));
 sky130_fd_sc_hd__dfxtp_2 _13003_ (.CLK(clk),
    .D(_01040_),
    .Q(\u_decod.branch_imm_q_o[16] ));
 sky130_fd_sc_hd__dfxtp_2 _13004_ (.CLK(clk),
    .D(_01041_),
    .Q(\u_decod.branch_imm_q_o[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clk),
    .D(_01042_),
    .Q(\u_decod.branch_imm_q_o[18] ));
 sky130_fd_sc_hd__dfxtp_2 _13006_ (.CLK(clk),
    .D(_01043_),
    .Q(\u_decod.branch_imm_q_o[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clk),
    .D(_01044_),
    .Q(\u_decod.branch_imm_q_o[20] ));
 sky130_fd_sc_hd__dfxtp_2 _13008_ (.CLK(clk),
    .D(_01045_),
    .Q(\u_decod.branch_imm_q_o[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clk),
    .D(_01046_),
    .Q(\u_decod.branch_imm_q_o[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clk),
    .D(_01047_),
    .Q(\u_decod.branch_imm_q_o[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13011_ (.CLK(clk),
    .D(_01048_),
    .Q(\u_decod.branch_imm_q_o[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13012_ (.CLK(clk),
    .D(_01049_),
    .Q(\u_decod.branch_imm_q_o[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clk),
    .D(_01050_),
    .Q(\u_decod.branch_imm_q_o[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clk),
    .D(_01051_),
    .Q(\u_decod.branch_imm_q_o[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clk),
    .D(_01052_),
    .Q(\u_decod.branch_imm_q_o[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clk),
    .D(_01053_),
    .Q(\u_decod.branch_imm_q_o[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clk),
    .D(_01054_),
    .Q(\u_decod.branch_imm_q_o[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clk),
    .D(_01055_),
    .Q(\u_decod.branch_imm_q_o[31] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_2955 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(icache_instr_i[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(icache_instr_i[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(icache_instr_i[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(icache_instr_i[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(icache_instr_i[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(icache_instr_i[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(icache_instr_i[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input8 (.A(icache_instr_i[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(icache_instr_i[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 input10 (.A(icache_instr_i[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(icache_instr_i[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(icache_instr_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(icache_instr_i[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(icache_instr_i[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(icache_instr_i[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(icache_instr_i[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(icache_instr_i[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(icache_instr_i[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(icache_instr_i[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(icache_instr_i[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(icache_instr_i[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(icache_instr_i[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(icache_instr_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(icache_instr_i[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(icache_instr_i[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(icache_instr_i[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(icache_instr_i[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(icache_instr_i[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(icache_instr_i[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(icache_instr_i[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(icache_instr_i[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(icache_instr_i[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(load_data_i[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(load_data_i[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(load_data_i[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(load_data_i[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(load_data_i[13]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(load_data_i[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(load_data_i[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(load_data_i[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(load_data_i[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(load_data_i[18]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(load_data_i[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(load_data_i[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(load_data_i[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(load_data_i[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(load_data_i[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 input48 (.A(load_data_i[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(load_data_i[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(load_data_i[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(load_data_i[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input52 (.A(load_data_i[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 input53 (.A(load_data_i[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(load_data_i[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(load_data_i[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(load_data_i[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(load_data_i[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(load_data_i[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(load_data_i[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(load_data_i[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(load_data_i[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(load_data_i[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(load_data_i[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(load_data_i[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(reset_adr_i[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(reset_adr_i[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(reset_adr_i[11]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(reset_adr_i[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(reset_adr_i[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(reset_adr_i[14]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(reset_adr_i[15]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(reset_adr_i[16]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(reset_adr_i[17]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(reset_adr_i[18]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(reset_adr_i[19]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(reset_adr_i[1]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(reset_adr_i[20]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(reset_adr_i[21]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(reset_adr_i[22]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(reset_adr_i[23]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(reset_adr_i[24]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(reset_adr_i[25]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(reset_adr_i[26]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(reset_adr_i[27]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(reset_adr_i[28]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(reset_adr_i[29]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(reset_adr_i[2]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(reset_adr_i[30]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(reset_adr_i[31]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input90 (.A(reset_adr_i[3]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(reset_adr_i[4]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(reset_adr_i[5]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(reset_adr_i[6]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(reset_adr_i[7]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(reset_adr_i[8]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(reset_adr_i[9]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(reset_n),
    .X(net97));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(access_size_o[0]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(access_size_o[1]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(access_size_o[2]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(adr_o[0]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(adr_o[10]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(adr_o[11]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(adr_o[12]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(adr_o[13]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(adr_o[14]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(adr_o[15]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(adr_o[16]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(adr_o[17]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(adr_o[18]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(adr_o[19]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(adr_o[1]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(adr_o[20]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(adr_o[21]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(adr_o[22]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(adr_o[23]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(adr_o[24]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(adr_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(adr_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(adr_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(adr_o[28]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(adr_o[29]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(adr_o[2]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(adr_o[30]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(adr_o[31]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(adr_o[3]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(adr_o[4]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(adr_o[5]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(adr_o[6]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(adr_o[7]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(adr_o[8]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(adr_o[9]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(adr_v_o));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(icache_adr_o[0]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(icache_adr_o[10]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(icache_adr_o[11]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(icache_adr_o[12]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(icache_adr_o[13]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(icache_adr_o[14]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(icache_adr_o[15]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(icache_adr_o[16]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(icache_adr_o[17]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(icache_adr_o[18]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(icache_adr_o[19]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(icache_adr_o[1]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(icache_adr_o[20]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(icache_adr_o[21]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(icache_adr_o[22]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(icache_adr_o[23]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(icache_adr_o[24]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(icache_adr_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(icache_adr_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(icache_adr_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(icache_adr_o[28]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(icache_adr_o[29]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(icache_adr_o[2]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(icache_adr_o[30]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(icache_adr_o[31]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(icache_adr_o[3]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(icache_adr_o[4]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(icache_adr_o[5]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(icache_adr_o[6]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(icache_adr_o[7]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(icache_adr_o[8]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(icache_adr_o[9]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(is_store_o));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(store_data_o[0]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(store_data_o[10]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(store_data_o[11]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(store_data_o[12]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(store_data_o[13]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(store_data_o[14]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(store_data_o[15]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(store_data_o[16]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(store_data_o[17]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(store_data_o[18]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(store_data_o[19]));
 sky130_fd_sc_hd__buf_2 output178 (.A(net178),
    .X(store_data_o[1]));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(store_data_o[20]));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net180),
    .X(store_data_o[21]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(store_data_o[22]));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(store_data_o[23]));
 sky130_fd_sc_hd__clkbuf_4 output183 (.A(net183),
    .X(store_data_o[24]));
 sky130_fd_sc_hd__clkbuf_4 output184 (.A(net184),
    .X(store_data_o[25]));
 sky130_fd_sc_hd__clkbuf_4 output185 (.A(net185),
    .X(store_data_o[26]));
 sky130_fd_sc_hd__clkbuf_4 output186 (.A(net186),
    .X(store_data_o[27]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(store_data_o[28]));
 sky130_fd_sc_hd__clkbuf_4 output188 (.A(net188),
    .X(store_data_o[29]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(store_data_o[2]));
 sky130_fd_sc_hd__clkbuf_4 output190 (.A(net190),
    .X(store_data_o[30]));
 sky130_fd_sc_hd__clkbuf_4 output191 (.A(net191),
    .X(store_data_o[31]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(store_data_o[3]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(store_data_o[4]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(store_data_o[5]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(store_data_o[6]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(store_data_o[7]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(store_data_o[8]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(store_data_o[9]));
 sky130_fd_sc_hd__clkbuf_2 max_cap199 (.A(_02085_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 max_cap200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 max_cap201 (.A(_01743_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net204),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_2 fanout204 (.A(net210),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_4 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_2 fanout207 (.A(net210),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(net210),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout210 (.A(net255),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(net220),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(net220),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net220),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net220),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(net219),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 fanout217 (.A(net219),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(net255),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_4 fanout221 (.A(net223),
    .X(net221));
 sky130_fd_sc_hd__buf_2 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(net255),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(net226),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(net255),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(net233),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net233),
    .X(net229));
 sky130_fd_sc_hd__buf_2 fanout230 (.A(net233),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_2 fanout233 (.A(net254),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(net238),
    .X(net234));
 sky130_fd_sc_hd__buf_2 fanout235 (.A(net238),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net254),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net254),
    .X(net239));
 sky130_fd_sc_hd__buf_2 fanout240 (.A(net254),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(net253),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 fanout242 (.A(net253),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net253),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net246),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 fanout246 (.A(net253),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 fanout248 (.A(net252),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(net252),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 fanout250 (.A(net252),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__buf_2 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 fanout255 (.A(net374),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net260),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(net260),
    .X(net258));
 sky130_fd_sc_hd__buf_2 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 fanout260 (.A(net270),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(net264),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 fanout264 (.A(net270),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 fanout266 (.A(net270),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_4 fanout267 (.A(net269),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_2 fanout270 (.A(net311),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(net274),
    .X(net271));
 sky130_fd_sc_hd__buf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(net311),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_2 fanout276 (.A(net311),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net279),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 fanout279 (.A(net311),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net283),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net283),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_2 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(net310),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 fanout284 (.A(net287),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_2 fanout285 (.A(net287),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_2 fanout287 (.A(net310),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net290),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(net310),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net293),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(net310),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net297),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_2 fanout295 (.A(net297),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(net310),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(net301),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_2 fanout299 (.A(net301),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_2 fanout301 (.A(net310),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 fanout302 (.A(net305),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(net305),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(net310),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(net309),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net374),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_4 fanout312 (.A(net318),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(net318),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(net318),
    .X(net314));
 sky130_fd_sc_hd__buf_2 fanout315 (.A(net318),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_4 fanout316 (.A(net318),
    .X(net316));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net334),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 fanout320 (.A(net334),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net334),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(net327),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 fanout324 (.A(net327),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_4 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net334),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_4 fanout328 (.A(net330),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_4 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net334),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net333),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 fanout334 (.A(net374),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_4 fanout335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__buf_2 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_2 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_4 fanout338 (.A(net374),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_4 fanout340 (.A(net348),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 fanout341 (.A(net348),
    .X(net341));
 sky130_fd_sc_hd__buf_2 fanout342 (.A(net343),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 fanout343 (.A(net348),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_4 fanout344 (.A(net348),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(net348),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(net348),
    .X(net346));
 sky130_fd_sc_hd__buf_2 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(net373),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 fanout349 (.A(net359),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_4 fanout351 (.A(net359),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 fanout352 (.A(net354),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_4 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_2 fanout354 (.A(net359),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 fanout355 (.A(net358),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net358),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_4 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__buf_2 fanout359 (.A(net373),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net367),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_4 fanout362 (.A(net367),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_2 fanout363 (.A(net367),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(net366),
    .X(net364));
 sky130_fd_sc_hd__buf_2 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_2 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_2 fanout367 (.A(net373),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(net373),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(net373),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_2 fanout372 (.A(net373),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_4 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_8 fanout374 (.A(net97),
    .X(net374));
endmodule
