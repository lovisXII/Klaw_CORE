* NGSPICE file created from core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt core VGND VPWR access_size_o[0] access_size_o[1] access_size_o[2] adr_o[0]
+ adr_o[10] adr_o[11] adr_o[12] adr_o[13] adr_o[14] adr_o[15] adr_o[16] adr_o[17]
+ adr_o[18] adr_o[19] adr_o[1] adr_o[20] adr_o[21] adr_o[22] adr_o[23] adr_o[24] adr_o[25]
+ adr_o[26] adr_o[27] adr_o[28] adr_o[29] adr_o[2] adr_o[30] adr_o[31] adr_o[3] adr_o[4]
+ adr_o[5] adr_o[6] adr_o[7] adr_o[8] adr_o[9] adr_v_o clk icache_adr_o[0] icache_adr_o[10]
+ icache_adr_o[11] icache_adr_o[12] icache_adr_o[13] icache_adr_o[14] icache_adr_o[15]
+ icache_adr_o[16] icache_adr_o[17] icache_adr_o[18] icache_adr_o[19] icache_adr_o[1]
+ icache_adr_o[20] icache_adr_o[21] icache_adr_o[22] icache_adr_o[23] icache_adr_o[24]
+ icache_adr_o[25] icache_adr_o[26] icache_adr_o[27] icache_adr_o[28] icache_adr_o[29]
+ icache_adr_o[2] icache_adr_o[30] icache_adr_o[31] icache_adr_o[3] icache_adr_o[4]
+ icache_adr_o[5] icache_adr_o[6] icache_adr_o[7] icache_adr_o[8] icache_adr_o[9]
+ icache_instr_i[0] icache_instr_i[10] icache_instr_i[11] icache_instr_i[12] icache_instr_i[13]
+ icache_instr_i[14] icache_instr_i[15] icache_instr_i[16] icache_instr_i[17] icache_instr_i[18]
+ icache_instr_i[19] icache_instr_i[1] icache_instr_i[20] icache_instr_i[21] icache_instr_i[22]
+ icache_instr_i[23] icache_instr_i[24] icache_instr_i[25] icache_instr_i[26] icache_instr_i[27]
+ icache_instr_i[28] icache_instr_i[29] icache_instr_i[2] icache_instr_i[30] icache_instr_i[31]
+ icache_instr_i[3] icache_instr_i[4] icache_instr_i[5] icache_instr_i[6] icache_instr_i[7]
+ icache_instr_i[8] icache_instr_i[9] is_store_o load_data_i[0] load_data_i[10] load_data_i[11]
+ load_data_i[12] load_data_i[13] load_data_i[14] load_data_i[15] load_data_i[16]
+ load_data_i[17] load_data_i[18] load_data_i[19] load_data_i[1] load_data_i[20] load_data_i[21]
+ load_data_i[22] load_data_i[23] load_data_i[24] load_data_i[25] load_data_i[26]
+ load_data_i[27] load_data_i[28] load_data_i[29] load_data_i[2] load_data_i[30] load_data_i[31]
+ load_data_i[3] load_data_i[4] load_data_i[5] load_data_i[6] load_data_i[7] load_data_i[8]
+ load_data_i[9] reset_adr_i[0] reset_adr_i[10] reset_adr_i[11] reset_adr_i[12] reset_adr_i[13]
+ reset_adr_i[14] reset_adr_i[15] reset_adr_i[16] reset_adr_i[17] reset_adr_i[18]
+ reset_adr_i[19] reset_adr_i[1] reset_adr_i[20] reset_adr_i[21] reset_adr_i[22] reset_adr_i[23]
+ reset_adr_i[24] reset_adr_i[25] reset_adr_i[26] reset_adr_i[27] reset_adr_i[28]
+ reset_adr_i[29] reset_adr_i[2] reset_adr_i[30] reset_adr_i[31] reset_adr_i[3] reset_adr_i[4]
+ reset_adr_i[5] reset_adr_i[6] reset_adr_i[7] reset_adr_i[8] reset_adr_i[9] reset_n
+ store_data_o[0] store_data_o[10] store_data_o[11] store_data_o[12] store_data_o[13]
+ store_data_o[14] store_data_o[15] store_data_o[16] store_data_o[17] store_data_o[18]
+ store_data_o[19] store_data_o[1] store_data_o[20] store_data_o[21] store_data_o[22]
+ store_data_o[23] store_data_o[24] store_data_o[25] store_data_o[26] store_data_o[27]
+ store_data_o[28] store_data_o[29] store_data_o[2] store_data_o[30] store_data_o[31]
+ store_data_o[3] store_data_o[4] store_data_o[5] store_data_o[6] store_data_o[7]
+ store_data_o[8] store_data_o[9]
XFILLER_0_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05903_ net510 _01118_ _01119_ net88 _01194_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__a221o_2
X_09671_ _04614_ VGND VGND VPWR VPWR _00133_ sky130_fd_sc_hd__clkbuf_1
X_06883_ _01305_ _01308_ _01341_ _01345_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__o31ai_2
X_08622_ u_rf.reg7_q\[21\] _03369_ _03370_ u_rf.reg25_q\[21\] _03804_ VGND VGND VPWR
+ VPWR _03805_ sky130_fd_sc_hd__a221o_1
X_05834_ _01104_ VGND VGND VPWR VPWR _01142_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_124_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08553_ u_rf.reg26_q\[18\] _03344_ _03282_ u_rf.reg10_q\[18\] _03738_ VGND VGND VPWR
+ VPWR _03739_ sky130_fd_sc_hd__a221o_1
X_05765_ _01086_ _01087_ VGND VGND VPWR VPWR _01088_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08484_ u_rf.reg4_q\[15\] _03265_ _03357_ u_rf.reg17_q\[15\] VGND VGND VPWR VPWR
+ _03673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07504_ _02619_ net47 _02446_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__a21bo_1
X_07435_ _01595_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07366_ u_rf.reg28_q\[19\] _01625_ _01631_ u_rf.reg17_q\[19\] _02597_ VGND VGND VPWR
+ VPWR _02598_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06317_ _01586_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_8
X_09105_ _04238_ _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07297_ _01381_ _01400_ _02443_ _01401_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__a31o_1
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06248_ _01517_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__inv_2
X_09036_ _01350_ _01345_ _01342_ _01347_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06179_ u_decod.rs2_data_q\[2\] VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09938_ _04768_ u_rf.reg7_q\[22\] _04764_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09869_ _04721_ VGND VGND VPWR VPWR _04722_ sky130_fd_sc_hd__buf_6
X_12880_ clknet_leaf_55_clk _00917_ net294 VGND VGND VPWR VPWR u_rf.reg28_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11900_ clknet_leaf_91_clk u_decod.rs2_data_nxt\[21\] net345 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[21\] sky130_fd_sc_hd__dfrtp_1
X_11831_ clknet_leaf_98_clk net19 net329 VGND VGND VPWR VPWR u_decod.dec0.funct7\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11762_ clknet_leaf_56_clk _00054_ net291 VGND VGND VPWR VPWR u_rf.reg1_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_509 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11693_ _05721_ VGND VGND VPWR VPWR _01048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10713_ u_rf.reg18_q\[12\] _04964_ _05199_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10644_ _05165_ VGND VGND VPWR VPWR _00555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10575_ u_rf.reg16_q\[11\] _04962_ _05127_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12314_ clknet_leaf_61_clk _00351_ net339 VGND VGND VPWR VPWR u_rf.reg10_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer7 _01113_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_1
X_12245_ clknet_leaf_45_clk _00282_ net300 VGND VGND VPWR VPWR u_rf.reg8_q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12176_ clknet_leaf_36_clk _00213_ net271 VGND VGND VPWR VPWR u_rf.reg6_q\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11127_ _05421_ VGND VGND VPWR VPWR _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11058_ _04751_ u_rf.reg23_q\[14\] _05380_ VGND VGND VPWR VPWR _05385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10009_ u_rf.reg8_q\[19\] _04467_ _04801_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_103_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07220_ _01422_ _02407_ _02458_ _01441_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__o211a_1
X_07151_ u_decod.rf_ff_res_data_i\[14\] _02358_ _02359_ _02390_ _02392_ VGND VGND
+ VPWR VPWR _02393_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06102_ u_decod.rs2_data_q\[22\] _01371_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07082_ _02309_ _02318_ _02325_ _01679_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06033_ _01301_ _01303_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07984_ u_decod.dec0.instr_i\[16\] VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09723_ _04641_ VGND VGND VPWR VPWR _00158_ sky130_fd_sc_hd__clkbuf_1
X_06935_ u_decod.pc_q_o\[11\] _02150_ _01484_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o21ai_1
X_09654_ _04604_ VGND VGND VPWR VPWR _00126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06866_ u_rf.reg31_q\[9\] _01614_ _01648_ u_rf.reg4_q\[9\] VGND VGND VPWR VPWR _02118_
+ sky130_fd_sc_hd__a22o_1
X_08605_ u_rf.reg28_q\[20\] _03556_ _03557_ u_rf.reg2_q\[20\] VGND VGND VPWR VPWR
+ _03789_ sky130_fd_sc_hd__a22o_1
X_05817_ u_decod.pc0_q_i\[9\] u_decod.pc0_q_i\[10\] _01124_ VGND VGND VPWR VPWR _01129_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_97_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ u_rf.reg0_q\[31\] _04492_ _04532_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__mux2_1
X_06797_ net63 _02047_ _02049_ net49 _02051_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08536_ u_rf.reg15_q\[17\] _03237_ _03302_ u_rf.reg24_q\[17\] _03722_ VGND VGND VPWR
+ VPWR _03723_ sky130_fd_sc_hd__a221o_1
X_05748_ u_decod.dec0.funct3\[0\] VGND VGND VPWR VPWR _01071_ sky130_fd_sc_hd__buf_2
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08467_ u_rf.reg28_q\[14\] _03242_ _03243_ u_rf.reg2_q\[14\] VGND VGND VPWR VPWR
+ _03657_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07418_ u_rf.reg27_q\[20\] _01671_ _01673_ u_rf.reg2_q\[20\] VGND VGND VPWR VPWR
+ _02648_ sky130_fd_sc_hd__a22o_1
X_08398_ u_rf.reg9_q\[11\] _03348_ _03349_ u_rf.reg20_q\[11\] VGND VGND VPWR VPWR
+ _03591_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07349_ _02536_ _02581_ _01424_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10360_ _04736_ u_rf.reg13_q\[7\] _05006_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09019_ _04163_ net406 VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__xor2_1
X_10291_ _04969_ VGND VGND VPWR VPWR _00398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12030_ clknet_leaf_113_clk u_decod.exe_ff_res_data_i\[10\] net328 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_57_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ clknet_leaf_106_clk _00969_ net320 VGND VGND VPWR VPWR u_rf.reg30_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12863_ clknet_leaf_133_clk _00900_ net231 VGND VGND VPWR VPWR u_rf.reg28_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12794_ clknet_leaf_93_clk _00831_ net340 VGND VGND VPWR VPWR u_rf.reg25_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11814_ clknet_leaf_95_clk net32 net331 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11745_ clknet_leaf_116_clk _00037_ net324 VGND VGND VPWR VPWR u_rf.reg1_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11676_ _05712_ VGND VGND VPWR VPWR _01040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10627_ _05156_ VGND VGND VPWR VPWR _00547_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10558_ u_rf.reg16_q\[3\] _04945_ _05116_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12228_ clknet_leaf_108_clk _00265_ net314 VGND VGND VPWR VPWR u_rf.reg8_q\[9\] sky130_fd_sc_hd__dfrtp_1
X_10489_ _05082_ VGND VGND VPWR VPWR _00483_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12159_ clknet_leaf_137_clk _00196_ net206 VGND VGND VPWR VPWR u_rf.reg6_q\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06720_ u_rf.reg1_q\[6\] _01586_ _01575_ u_rf.reg25_q\[6\] VGND VGND VPWR VPWR _01978_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06651_ _01479_ _01911_ _01441_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ u_rf.reg2_q\[6\] _04440_ _04428_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06582_ u_rf.reg30_q\[3\] _01579_ _01597_ u_rf.reg13_q\[3\] VGND VGND VPWR VPWR _01846_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08321_ u_rf.reg28_q\[7\] _03331_ _03333_ u_rf.reg2_q\[7\] VGND VGND VPWR VPWR _03518_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08252_ u_rf.reg27_q\[4\] _03319_ _03321_ u_rf.reg19_q\[4\] _03451_ VGND VGND VPWR
+ VPWR _03452_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07203_ _01357_ _01391_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
X_08183_ u_rf.reg1_q\[2\] _03310_ _03312_ u_rf.reg14_q\[2\] VGND VGND VPWR VPWR _03385_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07134_ _01598_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_136_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07065_ u_rf.reg16_q\[13\] _02307_ _01776_ u_rf.reg2_q\[13\] _02308_ VGND VGND VPWR
+ VPWR _02309_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06016_ _01277_ _01280_ _01283_ _01286_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__nand4_2
XFILLER_0_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_272 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07967_ u_decod.dec0.instr_i\[17\] u_decod.dec0.instr_i\[18\] VGND VGND VPWR VPWR
+ _03173_ sky130_fd_sc_hd__nor2_2
X_09706_ u_rf.reg4_q\[22\] _04474_ _04630_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06918_ u_rf.reg14_q\[10\] _01657_ _01669_ u_rf.reg27_q\[10\] VGND VGND VPWR VPWR
+ _02168_ sky130_fd_sc_hd__a22o_1
X_07898_ u_rf.reg30_q\[30\] _01581_ _02665_ u_rf.reg19_q\[30\] VGND VGND VPWR VPWR
+ _03108_ sky130_fd_sc_hd__a22o_1
X_09637_ u_rf.reg3_q\[22\] _04474_ _04593_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__mux2_1
X_06849_ _01995_ _02101_ _01315_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__mux2_1
X_09568_ _04558_ VGND VGND VPWR VPWR _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ u_rf.reg0_q\[16\] _03420_ _03329_ u_rf.reg12_q\[16\] _03706_ VGND VGND VPWR
+ VPWR _03707_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_156_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _04521_ VGND VGND VPWR VPWR _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11530_ _04747_ u_rf.reg30_q\[12\] _05632_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_355 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11461_ _05598_ VGND VGND VPWR VPWR _00939_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10412_ _04423_ _04425_ _04936_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__or3_4
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11392_ u_rf.reg28_q\[11\] u_decod.rf_ff_res_data_i\[11\] _05560_ VGND VGND VPWR
+ VPWR _05562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10343_ _05004_ VGND VGND VPWR VPWR _00415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10274_ u_rf.reg12_q\[9\] _04957_ _04939_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__mux2_1
X_12013_ clknet_leaf_76_clk u_exe.bu_pc_res\[26\] net369 VGND VGND VPWR VPWR u_exe.pc_data_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12915_ clknet_leaf_68_clk _00952_ net351 VGND VGND VPWR VPWR u_rf.reg29_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ clknet_leaf_7_clk _00883_ net218 VGND VGND VPWR VPWR u_rf.reg27_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_732 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12777_ clknet_leaf_20_clk _00814_ net283 VGND VGND VPWR VPWR u_rf.reg25_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11728_ clknet_leaf_35_clk _00020_ net271 VGND VGND VPWR VPWR u_rf.reg2_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11659_ _05693_ u_decod.branch_imm_q_o\[8\] VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08870_ _04035_ _04036_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07821_ u_rf.reg31_q\[28\] _01777_ _02385_ u_rf.reg20_q\[28\] _03034_ VGND VGND VPWR
+ VPWR _03035_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07752_ _01746_ _02966_ _02968_ _01260_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__a22o_1
X_07683_ _02893_ _02902_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__or2_1
X_06703_ u_decod.pc_q_o\[6\] _01917_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__or2_1
X_09422_ u_decod.rf_ff_res_data_i\[23\] VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__buf_2
X_06634_ _01075_ _01740_ _01741_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09353_ _04429_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06565_ _01810_ _01822_ _01829_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__or3_1
XFILLER_0_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08304_ u_rf.reg8_q\[7\] _03407_ _03408_ u_rf.reg29_q\[7\] _03500_ VGND VGND VPWR
+ VPWR _03501_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06496_ u_decod.instr_operation_q\[1\] _01259_ VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__nand2_4
XFILLER_0_7_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09284_ _04385_ u_decod.rs2_data_q\[5\] _04386_ VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08235_ u_rf.reg4_q\[4\] _03265_ _03267_ u_rf.reg17_q\[4\] VGND VGND VPWR VPWR _03435_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08166_ _03229_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_151_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07117_ _01680_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08097_ _03300_ VGND VGND VPWR VPWR _03301_ sky130_fd_sc_hd__buf_8
X_07048_ u_decod.rs1_data_q\[13\] _01454_ _01685_ _02136_ VGND VGND VPWR VPWR _02293_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_54_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08999_ u_decod.rs1_data_q\[27\] u_decod.branch_imm_q_o\[27\] VGND VGND VPWR VPWR
+ _04147_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10961_ u_rf.reg22_q\[0\] _04935_ _05333_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12700_ clknet_leaf_129_clk _00737_ net234 VGND VGND VPWR VPWR u_rf.reg23_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12631_ clknet_leaf_70_clk _00668_ net352 VGND VGND VPWR VPWR u_rf.reg20_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_10892_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__buf_6
XFILLER_0_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12562_ clknet_leaf_40_clk _00599_ net278 VGND VGND VPWR VPWR u_rf.reg18_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12493_ clknet_leaf_5_clk _00530_ net217 VGND VGND VPWR VPWR u_rf.reg16_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_11513_ _04730_ u_rf.reg30_q\[4\] _05621_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11444_ _05589_ VGND VGND VPWR VPWR _00931_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11375_ u_rf.reg28_q\[3\] net491 _05549_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10326_ u_decod.rf_ff_res_data_i\[26\] VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10257_ _04946_ VGND VGND VPWR VPWR _00387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10188_ _04734_ u_rf.reg11_q\[6\] _04900_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_58 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12829_ clknet_leaf_13_clk _00866_ net244 VGND VGND VPWR VPWR u_rf.reg27_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06350_ _01572_ _01514_ _01573_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__and3_2
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06281_ _01522_ u_decod.dec0.instr_i\[23\] VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__nor2_2
XFILLER_0_16_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08020_ u_rf.reg4_q\[31\] _03224_ _03225_ u_rf.reg17_q\[31\] VGND VGND VPWR VPWR
+ _03226_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09971_ _04791_ VGND VGND VPWR VPWR _00256_ sky130_fd_sc_hd__clkbuf_1
X_08922_ _04074_ _04077_ _04073_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_110_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08853_ _03998_ _04022_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__nor2_1
XFILLER_0_34_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08784_ u_rf.reg28_q\[29\] _03556_ _03356_ u_rf.reg4_q\[29\] _03958_ VGND VGND VPWR
+ VPWR _03959_ sky130_fd_sc_hd__a221o_1
X_07804_ _02334_ _02998_ _02999_ _03018_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__o31a_1
XFILLER_0_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05996_ u_decod.rs1_data_q\[31\] VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__buf_4
X_07735_ _01528_ _02840_ _02861_ _02906_ VGND VGND VPWR VPWR _02953_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_28_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07666_ u_rf.reg6_q\[25\] _01556_ _01630_ u_rf.reg17_q\[25\] _02885_ VGND VGND VPWR
+ VPWR _02886_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09405_ _04464_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07597_ _01280_ VGND VGND VPWR VPWR _02820_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06617_ u_rf.reg31_q\[4\] _01615_ _01649_ u_rf.reg4_q\[4\] VGND VGND VPWR VPWR _01879_
+ sky130_fd_sc_hd__a22o_1
X_09336_ _04409_ u_decod.rs2_data_q\[29\] _04410_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06548_ _01812_ _01312_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__nor2_1
X_09267_ _04372_ _04374_ VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06479_ _01506_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08218_ _03412_ _03414_ _03416_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__or4_1
X_09198_ _04307_ _04314_ _04312_ _04319_ _04311_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a311o_1
XFILLER_0_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08149_ _03222_ VGND VGND VPWR VPWR _03352_ sky130_fd_sc_hd__buf_6
XFILLER_0_114_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11160_ _05438_ VGND VGND VPWR VPWR _00798_ sky130_fd_sc_hd__clkbuf_1
X_11091_ _04784_ u_rf.reg23_q\[30\] _05368_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__mux2_1
X_10111_ u_rf.reg10_q\[2\] _04432_ _04863_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__mux2_1
X_10042_ _04829_ VGND VGND VPWR VPWR _00289_ sky130_fd_sc_hd__clkbuf_1
Xhold74 u_decod.pc0_q_i\[11\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 u_decod.exe_ff_rd_adr_q_i\[1\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold85 u_decod.pc0_q_i\[12\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 u_decod.pc0_q_i\[10\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ clknet_leaf_84_clk u_exe.bu_pc_res\[6\] net364 VGND VGND VPWR VPWR u_exe.pc_data_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10944_ _05324_ VGND VGND VPWR VPWR _00696_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10875_ _05287_ VGND VGND VPWR VPWR _00664_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12614_ clknet_leaf_0_clk _00651_ net203 VGND VGND VPWR VPWR u_rf.reg20_q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12545_ clknet_leaf_95_clk _00582_ net325 VGND VGND VPWR VPWR u_rf.reg18_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_132_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_132_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12476_ clknet_leaf_127_clk _00513_ net237 VGND VGND VPWR VPWR u_rf.reg16_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11427_ u_rf.reg28_q\[28\] u_decod.rf_ff_res_data_i\[28\] _05571_ VGND VGND VPWR
+ VPWR _05580_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 _01554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11358_ _05543_ VGND VGND VPWR VPWR _00891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10309_ u_rf.reg12_q\[20\] _04980_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11289_ u_rf.reg26_q\[27\] u_decod.rf_ff_res_data_i\[27\] _05499_ VGND VGND VPWR
+ VPWR _05507_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05850_ _01153_ _01144_ _01154_ VGND VGND VPWR VPWR _01155_ sky130_fd_sc_hd__and3b_1
XFILLER_0_83_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer17 u_decod.pc0_q_i\[2\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07520_ u_rf.reg3_q\[22\] _02363_ _02697_ u_rf.reg4_q\[22\] _02745_ VGND VGND VPWR
+ VPWR _02746_ sky130_fd_sc_hd__a221o_1
Xrebuffer28 net403 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
X_05781_ u_decod.pc0_q_i\[0\] _01099_ _01101_ net65 _01102_ VGND VGND VPWR VPWR net134
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_79 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07451_ _02493_ _02679_ _01472_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07382_ _02603_ _02613_ _01680_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__o21a_2
XFILLER_0_18_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06402_ _01513_ _01515_ _01553_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__and3_2
X_09121_ _04253_ _04248_ _04245_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__o21a_1
XFILLER_0_85_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06333_ u_rf.reg18_q\[0\] _01592_ _01595_ u_rf.reg19_q\[0\] _01602_ VGND VGND VPWR
+ VPWR _01603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_123_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_123_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_98_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09052_ u_decod.instr_operation_q\[5\] VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__inv_2
X_06264_ u_decod.rf_ff_rd_adr_q_i\[0\] VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08003_ u_decod.dec0.instr_i\[15\] u_decod.dec0.instr_i\[16\] VGND VGND VPWR VPWR
+ _03209_ sky130_fd_sc_hd__and2_2
X_06195_ _01461_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_386 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09954_ _04779_ VGND VGND VPWR VPWR _00251_ sky130_fd_sc_hd__clkbuf_1
X_08905_ u_decod.rs1_data_q\[13\] u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR
+ _04067_ sky130_fd_sc_hd__nor2_1
X_09885_ _04732_ u_rf.reg7_q\[5\] _04722_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_146_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ u_decod.rs1_data_q\[2\] u_decod.branch_imm_q_o\[2\] VGND VGND VPWR VPWR _04008_
+ sky130_fd_sc_hd__or2_1
X_08767_ u_rf.reg30_q\[28\] _03281_ _03283_ u_rf.reg10_q\[28\] _03942_ VGND VGND VPWR
+ VPWR _03943_ sky130_fd_sc_hd__a221o_1
X_05979_ _01234_ _01253_ VGND VGND VPWR VPWR _01254_ sky130_fd_sc_hd__and2_1
X_07718_ u_rf.reg29_q\[26\] _01780_ _02697_ u_rf.reg4_q\[26\] _02935_ VGND VGND VPWR
+ VPWR _02936_ sky130_fd_sc_hd__a221o_1
X_08698_ u_rf.reg18_q\[25\] _03262_ _03263_ u_rf.reg23_q\[25\] _03876_ VGND VGND VPWR
+ VPWR _03877_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07649_ _02786_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__inv_2
X_10660_ _05173_ VGND VGND VPWR VPWR _00563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09319_ _04407_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_149_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10591_ u_rf.reg16_q\[19\] _04978_ _05127_ VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_114_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_114_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_11_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12330_ clknet_leaf_30_clk _00367_ net262 VGND VGND VPWR VPWR u_rf.reg11_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ clknet_leaf_125_clk _00298_ net239 VGND VGND VPWR VPWR u_rf.reg9_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11212_ _05466_ VGND VGND VPWR VPWR _00822_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12192_ clknet_leaf_117_clk _00229_ net324 VGND VGND VPWR VPWR u_rf.reg7_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_11143_ u_rf.reg24_q\[22\] _04985_ _05427_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__mux2_1
X_11074_ _05393_ VGND VGND VPWR VPWR _00757_ sky130_fd_sc_hd__clkbuf_1
X_10025_ _04819_ VGND VGND VPWR VPWR _00282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11976_ clknet_leaf_75_clk net455 net368 VGND VGND VPWR VPWR u_decod.pc_q_o\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10927_ _05315_ VGND VGND VPWR VPWR _00688_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_510 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10858_ _05278_ VGND VGND VPWR VPWR _00656_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_105_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_105_clk sky130_fd_sc_hd__clkbuf_16
X_10789_ net521 _04972_ _05235_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12528_ clknet_leaf_31_clk _00565_ net263 VGND VGND VPWR VPWR u_rf.reg17_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12459_ clknet_leaf_136_clk _00496_ net207 VGND VGND VPWR VPWR u_rf.reg15_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout309 net310 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06951_ _01424_ _02198_ _02199_ _01506_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__o211a_1
X_05902_ _01192_ _01098_ _01193_ VGND VGND VPWR VPWR _01194_ sky130_fd_sc_hd__and3b_1
X_09670_ u_rf.reg4_q\[5\] _04438_ _04608_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__mux2_1
X_08621_ u_rf.reg1_q\[21\] _03310_ _03312_ u_rf.reg14_q\[21\] VGND VGND VPWR VPWR
+ _03804_ sky130_fd_sc_hd__a22o_1
X_06882_ _02132_ _02133_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[9\] sky130_fd_sc_hd__xnor2_1
X_05833_ net507 _01105_ _01132_ net69 _01141_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_124_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ u_rf.reg28_q\[18\] _03330_ _03217_ u_rf.reg29_q\[18\] VGND VGND VPWR VPWR
+ _03738_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05764_ u_decod.dec0.instr_i\[6\] u_decod.dec0.instr_i\[5\] VGND VGND VPWR VPWR _01087_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ u_rf.reg8_q\[15\] _03407_ _03408_ u_rf.reg29_q\[15\] _03671_ VGND VGND VPWR
+ VPWR _03672_ sky130_fd_sc_hd__a221o_1
X_07503_ _02723_ _02682_ _02729_ _01443_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07434_ _01569_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07365_ u_rf.reg31_q\[19\] _01615_ _01622_ u_rf.reg24_q\[19\] VGND VGND VPWR VPWR
+ _02597_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09104_ u_decod.pc_q_o\[7\] u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _04239_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07296_ _02530_ _02531_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[17\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06316_ _01585_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__buf_6
X_09035_ _01314_ _01426_ _01766_ _01813_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06247_ u_decod.dec0.instr_i\[6\] u_decod.dec0.instr_i\[4\] _01225_ _01516_ VGND
+ VGND VPWR VPWR _01517_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06178_ u_decod.rs1_data_q\[7\] _01289_ _01367_ _01267_ _01444_ _01447_ VGND VGND
+ VPWR VPWR _01449_ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09937_ u_decod.rf_ff_res_data_i\[22\] VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09868_ _04720_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__clkbuf_4
X_08819_ u_rf.reg7_q\[30\] _03314_ _03315_ u_rf.reg25_q\[30\] _03992_ VGND VGND VPWR
+ VPWR _03993_ sky130_fd_sc_hd__a221o_1
X_09799_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__buf_8
XFILLER_0_96_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11830_ clknet_leaf_98_clk net18 net329 VGND VGND VPWR VPWR u_decod.dec0.funct7\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_157_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11761_ clknet_leaf_35_clk _00053_ net271 VGND VGND VPWR VPWR u_rf.reg1_q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10712_ _05201_ VGND VGND VPWR VPWR _00587_ sky130_fd_sc_hd__clkbuf_1
X_11692_ u_decod.branch_imm_q_o\[24\] _02841_ _05717_ VGND VGND VPWR VPWR _05721_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10643_ u_rf.reg17_q\[11\] _04962_ _05163_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10574_ _05128_ VGND VGND VPWR VPWR _00522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12313_ clknet_leaf_63_clk _00350_ net342 VGND VGND VPWR VPWR u_rf.reg10_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer8 _01113_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12244_ clknet_leaf_33_clk _00281_ net269 VGND VGND VPWR VPWR u_rf.reg8_q\[25\] sky130_fd_sc_hd__dfrtp_1
X_12175_ clknet_leaf_35_clk _00212_ net272 VGND VGND VPWR VPWR u_rf.reg6_q\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11126_ u_rf.reg24_q\[14\] _04968_ _05416_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11057_ _05384_ VGND VGND VPWR VPWR _00749_ sky130_fd_sc_hd__clkbuf_1
X_10008_ _04810_ VGND VGND VPWR VPWR _00274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11959_ clknet_leaf_101_clk net474 net374 VGND VGND VPWR VPWR u_decod.pc_q_o\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07150_ _02305_ _02391_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06101_ u_decod.rs2_data_q\[22\] _01371_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_95_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07081_ _02320_ _02322_ _02324_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06032_ u_decod.rs2_data_q\[10\] _01302_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ u_rf.reg4_q\[30\] _04490_ _04607_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__mux2_1
X_07983_ _01542_ u_decod.dec0.instr_i\[16\] _03181_ _01531_ VGND VGND VPWR VPWR _03189_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06934_ net35 _02047_ _02049_ net52 _02051_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__a221o_1
X_09653_ u_rf.reg3_q\[30\] _04490_ _04570_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__mux2_1
X_06865_ u_rf.reg29_q\[9\] _01626_ _01637_ u_rf.reg21_q\[9\] _02116_ VGND VGND VPWR
+ VPWR _02117_ sky130_fd_sc_hd__a221o_1
X_08604_ u_rf.reg27_q\[20\] _03319_ _03321_ u_rf.reg19_q\[20\] _03787_ VGND VGND VPWR
+ VPWR _03788_ sky130_fd_sc_hd__a221o_1
X_09584_ _04566_ VGND VGND VPWR VPWR _00094_ sky130_fd_sc_hd__clkbuf_1
X_05816_ net467 _01105_ _01101_ net96 _01128_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__a221o_1
XFILLER_0_96_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08535_ u_rf.reg6_q\[17\] _03235_ _03236_ u_rf.reg13_q\[17\] VGND VGND VPWR VPWR
+ _03722_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06796_ _02050_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_46_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05747_ net466 _01070_ VGND VGND VPWR VPWR u_decod.dec0.jalr sky130_fd_sc_hd__nor2_1
X_08466_ _03651_ _03653_ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__or3_1
X_07417_ u_decod.dec0.instr_i\[20\] _01206_ _02646_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08397_ u_rf.reg18_q\[11\] _03353_ _03355_ u_rf.reg23_q\[11\] _03589_ VGND VGND VPWR
+ VPWR _03590_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07348_ _02494_ _02580_ _01757_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07279_ u_rf.reg31_q\[17\] _01615_ _01658_ u_rf.reg14_q\[17\] _02514_ VGND VGND VPWR
+ VPWR _02515_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09018_ _04156_ _04157_ _04158_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__o21ai_2
X_10290_ u_rf.reg12_q\[14\] _04968_ _04960_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_57_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ clknet_leaf_106_clk _00968_ net319 VGND VGND VPWR VPWR u_rf.reg30_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12862_ clknet_leaf_123_clk _00899_ net241 VGND VGND VPWR VPWR u_rf.reg28_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11813_ clknet_leaf_95_clk net31 net331 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ clknet_leaf_64_clk _00830_ net346 VGND VGND VPWR VPWR u_rf.reg25_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11744_ clknet_leaf_131_clk _00036_ net227 VGND VGND VPWR VPWR u_rf.reg1_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11675_ u_decod.branch_imm_q_o\[16\] _02465_ _05696_ VGND VGND VPWR VPWR _05712_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10626_ u_rf.reg17_q\[3\] _04945_ _05152_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10557_ _05119_ VGND VGND VPWR VPWR _00514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10488_ _04728_ u_rf.reg15_q\[3\] _05078_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__mux2_1
X_12227_ clknet_leaf_108_clk _00264_ net314 VGND VGND VPWR VPWR u_rf.reg8_q\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12158_ clknet_leaf_134_clk _00195_ net209 VGND VGND VPWR VPWR u_rf.reg6_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_12089_ clknet_leaf_57_clk _00126_ net291 VGND VGND VPWR VPWR u_rf.reg3_q\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11109_ u_rf.reg24_q\[6\] _04951_ _05405_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_218 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06650_ _01807_ _01910_ _01688_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06581_ u_rf.reg23_q\[3\] _01613_ _01638_ u_rf.reg21_q\[3\] _01844_ VGND VGND VPWR
+ VPWR _01845_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08320_ u_rf.reg27_q\[7\] _03319_ _03321_ u_rf.reg19_q\[7\] _03516_ VGND VGND VPWR
+ VPWR _03517_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08251_ u_rf.reg16_q\[4\] _03450_ _03325_ u_rf.reg5_q\[4\] VGND VGND VPWR VPWR _03451_
+ sky130_fd_sc_hd__a22o_1
X_07202_ _02440_ _02441_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[15\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08182_ u_rf.reg0_q\[2\] _03176_ _03329_ u_rf.reg12_q\[2\] _03383_ VGND VGND VPWR
+ VPWR _03384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_389 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07133_ _01584_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_119_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_754 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07064_ u_rf.reg1_q\[13\] _01587_ _01667_ u_rf.reg8_q\[13\] VGND VGND VPWR VPWR _02308_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06015_ _01284_ _01285_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07966_ u_decod.dec0.instr_i\[15\] u_decod.dec0.instr_i\[16\] VGND VGND VPWR VPWR
+ _03172_ sky130_fd_sc_hd__nor2_2
X_09705_ _04632_ VGND VGND VPWR VPWR _00149_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06917_ u_rf.reg12_q\[10\] _01607_ _01672_ u_rf.reg2_q\[10\] _02166_ VGND VGND VPWR
+ VPWR _02167_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09636_ _04595_ VGND VGND VPWR VPWR _00117_ sky130_fd_sc_hd__clkbuf_1
X_07897_ u_rf.reg13_q\[30\] _02376_ _02386_ u_rf.reg27_q\[30\] _03106_ VGND VGND VPWR
+ VPWR _03107_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_94_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
X_06848_ _01909_ _02100_ _01450_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09567_ u_rf.reg0_q\[22\] _04474_ _04555_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06779_ _01772_ u_decod.exe_ff_res_data_i\[7\] _02034_ VGND VGND VPWR VPWR _02035_
+ sky130_fd_sc_hd__a21o_1
X_09498_ u_rf.reg1_q\[22\] _04474_ _04518_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ u_rf.reg28_q\[16\] _03556_ _03557_ u_rf.reg2_q\[16\] VGND VGND VPWR VPWR
+ _03706_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08449_ u_rf.reg24_q\[13\] _03238_ _03306_ u_rf.reg13_q\[13\] VGND VGND VPWR VPWR
+ _03640_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_671 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11460_ _04745_ u_rf.reg29_q\[11\] _05596_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__mux2_1
X_10411_ _05040_ VGND VGND VPWR VPWR _00447_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ _05561_ VGND VGND VPWR VPWR _00906_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10342_ u_rf.reg12_q\[31\] _05003_ _04938_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12012_ clknet_leaf_76_clk u_exe.bu_pc_res\[25\] net368 VGND VGND VPWR VPWR u_exe.pc_data_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10273_ u_decod.rf_ff_res_data_i\[9\] VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_131_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_85_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
X_12914_ clknet_leaf_39_clk _00951_ net279 VGND VGND VPWR VPWR u_rf.reg29_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12845_ clknet_leaf_11_clk _00882_ net224 VGND VGND VPWR VPWR u_rf.reg27_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_914 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12776_ clknet_leaf_17_clk _00813_ net289 VGND VGND VPWR VPWR u_rf.reg25_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11727_ clknet_leaf_6_clk _00019_ net216 VGND VGND VPWR VPWR u_rf.reg2_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_140_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11658_ u_decod.dec0.funct7\[2\] _05700_ _02644_ _05703_ VGND VGND VPWR VPWR _01031_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_490 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10609_ _05146_ VGND VGND VPWR VPWR _00539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_663 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11589_ _04738_ u_rf.reg31_q\[8\] _05657_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07820_ u_rf.reg1_q\[28\] _02604_ _02376_ u_rf.reg13_q\[28\] VGND VGND VPWR VPWR
+ _03034_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07751_ _01430_ _01282_ _01283_ u_decod.instr_operation_q\[3\] _02967_ VGND VGND
+ VPWR VPWR _02968_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_76_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06702_ u_decod.rs2_data_q\[6\] u_decod.rs1_data_q\[6\] VGND VGND VPWR VPWR _01961_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_126_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07682_ _02895_ _02897_ _02899_ _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09421_ _04475_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__clkbuf_1
X_06633_ _01713_ u_decod.exe_ff_res_data_i\[4\] _01894_ VGND VGND VPWR VPWR _01895_
+ sky130_fd_sc_hd__a21o_1
X_09352_ u_rf.reg2_q\[0\] _04421_ _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__mux2_1
X_06564_ _01506_ _01826_ _01828_ _01059_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08303_ u_rf.reg22_q\[7\] _03409_ _03410_ u_rf.reg3_q\[7\] VGND VGND VPWR VPWR _03500_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_138_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06495_ net55 _01487_ _01488_ net42 _01761_ VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09283_ _04388_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_1
XFILLER_0_145_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08234_ net389 _03259_ _03434_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[3\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08165_ u_rf.reg27_q\[1\] _03365_ _03366_ u_rf.reg19_q\[1\] _03367_ VGND VGND VPWR
+ VPWR _03368_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07116_ _01550_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__buf_4
XFILLER_0_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08096_ _03237_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__buf_6
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07047_ _02001_ _02197_ _01458_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08998_ _04101_ _04146_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_67_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
X_07949_ u_rf.reg7_q\[31\] _01562_ _02363_ u_rf.reg3_q\[31\] VGND VGND VPWR VPWR _03157_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10960_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__buf_6
X_09619_ _04586_ VGND VGND VPWR VPWR _00109_ sky130_fd_sc_hd__clkbuf_1
X_10891_ _04644_ _04645_ _05295_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__and3_2
X_12630_ clknet_leaf_51_clk _00667_ net308 VGND VGND VPWR VPWR u_rf.reg20_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12561_ clknet_leaf_56_clk _00598_ net291 VGND VGND VPWR VPWR u_rf.reg18_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12492_ clknet_leaf_25_clk _00529_ net265 VGND VGND VPWR VPWR u_rf.reg16_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11512_ _05625_ VGND VGND VPWR VPWR _00963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11443_ _04728_ u_rf.reg29_q\[3\] _05585_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11374_ _05552_ VGND VGND VPWR VPWR _00898_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10325_ _04992_ VGND VGND VPWR VPWR _00409_ sky130_fd_sc_hd__clkbuf_1
X_10256_ u_rf.reg12_q\[3\] _04945_ _04939_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10187_ _04906_ VGND VGND VPWR VPWR _00357_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_58_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_85_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12828_ clknet_leaf_128_clk _00865_ net237 VGND VGND VPWR VPWR u_rf.reg27_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12759_ clknet_leaf_70_clk _00796_ net352 VGND VGND VPWR VPWR u_rf.reg24_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06280_ _01549_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__buf_4
XFILLER_0_142_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09970_ u_rf.reg8_q\[0\] _04421_ _04790_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__mux2_1
X_08921_ _04079_ _04080_ VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__nor2_1
X_08852_ _04020_ _04021_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07803_ _01260_ _03006_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_49_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ u_rf.reg21_q\[29\] _03206_ _03211_ u_rf.reg11_q\[29\] VGND VGND VPWR VPWR
+ _03958_ sky130_fd_sc_hd__a22o_1
X_05995_ _01264_ _01265_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07734_ _01528_ _02929_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07665_ u_rf.reg13_q\[25\] _01597_ _01656_ u_rf.reg10_q\[25\] VGND VGND VPWR VPWR
+ _02885_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09404_ u_rf.reg2_q\[17\] _04463_ _04449_ VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06616_ u_rf.reg13_q\[4\] _01597_ _01592_ u_rf.reg18_q\[4\] _01877_ VGND VGND VPWR
+ VPWR _01878_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07596_ _02818_ _01405_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09335_ _04416_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_1
X_06547_ u_decod.rs1_data_q\[3\] _01468_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__and2_1
X_09266_ u_decod.pc_q_o\[30\] u_decod.branch_imm_q_o\[30\] VGND VGND VPWR VPWR _04378_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06478_ _01737_ _01745_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[1\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08217_ u_rf.reg30_q\[3\] _03341_ _03342_ u_rf.reg10_q\[3\] _03417_ VGND VGND VPWR
+ VPWR _03418_ sky130_fd_sc_hd__a221o_1
X_09197_ _04317_ _04318_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08148_ u_rf.reg31_q\[1\] _03290_ _03292_ u_rf.reg11_q\[1\] _03350_ VGND VGND VPWR
+ VPWR _03351_ sky130_fd_sc_hd__a221o_1
X_08079_ _03282_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__buf_8
XFILLER_0_113_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11090_ _05401_ VGND VGND VPWR VPWR _00765_ sky130_fd_sc_hd__clkbuf_1
X_10110_ _04865_ VGND VGND VPWR VPWR _00321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10041_ u_rf.reg9_q\[1\] _04430_ _04827_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__mux2_1
Xhold64 u_decod.pc0_q_i\[22\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 u_exe.pc_data_q\[14\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ clknet_leaf_87_clk u_exe.bu_pc_res\[5\] net362 VGND VGND VPWR VPWR u_exe.pc_data_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold75 u_decod.exe_ff_rd_adr_q_i\[2\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 u_decod.rf_ff_res_data_i\[9\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ u_rf.reg21_q\[24\] _04989_ _05319_ VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ u_rf.reg20_q\[24\] _04989_ _05282_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12613_ clknet_leaf_125_clk _00650_ net316 VGND VGND VPWR VPWR u_rf.reg20_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ clknet_leaf_116_clk _00581_ net323 VGND VGND VPWR VPWR u_rf.reg18_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12475_ clknet_leaf_10_clk _00512_ net224 VGND VGND VPWR VPWR u_rf.reg16_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11426_ _05579_ VGND VGND VPWR VPWR _00923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_6 _01561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11357_ _04778_ u_rf.reg27_q\[27\] _05535_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10308_ _04938_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__buf_6
XFILLER_0_67_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11288_ _05506_ VGND VGND VPWR VPWR _00858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _04933_ VGND VGND VPWR VPWR _00382_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer18 net410 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
X_05780_ u_decod.flush_v net360 net492 VGND VGND VPWR VPWR _01102_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer29 net404 VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07450_ _01468_ _02287_ _01498_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__o21a_1
XFILLER_0_146_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07381_ _02606_ _02608_ _02610_ _02612_ VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__or4_1
X_06401_ _01670_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09120_ _04246_ VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__inv_2
X_06332_ u_rf.reg13_q\[0\] _01598_ _01601_ u_rf.reg15_q\[0\] VGND VGND VPWR VPWR _01602_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09051_ _04190_ _04193_ _01485_ VGND VGND VPWR VPWR u_exe.branch_v sky130_fd_sc_hd__o21a_1
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08002_ u_rf.reg30_q\[31\] _03200_ _03202_ u_rf.reg10_q\[31\] _03207_ VGND VGND VPWR
+ VPWR _03208_ sky130_fd_sc_hd__a221o_1
X_06263_ u_decod.rf_ff_rd_adr_q_i\[0\] _01520_ u_decod.dec0.instr_i\[22\] _01532_
+ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06194_ _01462_ _01463_ _01464_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09953_ _04778_ u_rf.reg7_q\[27\] _04764_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08904_ _04042_ _04066_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__nor2_2
X_09884_ u_decod.rf_ff_res_data_i\[5\] VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_146_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _04005_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08766_ u_rf.reg26_q\[28\] _03284_ _03286_ u_rf.reg21_q\[28\] VGND VGND VPWR VPWR
+ _03942_ sky130_fd_sc_hd__a22o_1
X_07717_ u_rf.reg12_q\[26\] _01609_ _02368_ u_rf.reg26_q\[26\] VGND VGND VPWR VPWR
+ _02935_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05978_ _01074_ _01221_ _01252_ _01095_ VGND VGND VPWR VPWR _01253_ sky130_fd_sc_hd__a31o_1
X_08697_ u_rf.reg4_q\[25\] _03264_ _03266_ u_rf.reg17_q\[25\] VGND VGND VPWR VPWR
+ _03876_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07648_ u_decod.pc_q_o\[25\] _02816_ _01485_ VGND VGND VPWR VPWR _02869_ sky130_fd_sc_hd__o21ai_1
X_07579_ u_rf.reg5_q\[23\] _02664_ _02665_ u_rf.reg19_q\[23\] _02802_ VGND VGND VPWR
+ VPWR _02803_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09318_ _04397_ u_decod.rs2_data_q\[21\] _04398_ VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_62_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10590_ _05136_ VGND VGND VPWR VPWR _00530_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09249_ _04340_ _04345_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12260_ clknet_leaf_108_clk _00297_ net312 VGND VGND VPWR VPWR u_rf.reg9_q\[9\] sky130_fd_sc_hd__dfrtp_1
X_11211_ u_rf.reg25_q\[22\] _04985_ _05463_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__mux2_1
X_12191_ clknet_leaf_132_clk _00228_ net228 VGND VGND VPWR VPWR u_rf.reg7_q\[4\] sky130_fd_sc_hd__dfrtp_1
X_11142_ _05429_ VGND VGND VPWR VPWR _00789_ sky130_fd_sc_hd__clkbuf_1
X_11073_ _04766_ u_rf.reg23_q\[21\] _05391_ VGND VGND VPWR VPWR _05393_ sky130_fd_sc_hd__mux2_1
Xoutput98 net98 VGND VGND VPWR VPWR access_size_o[0] sky130_fd_sc_hd__buf_2
X_10024_ u_rf.reg8_q\[26\] _04482_ _04812_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__mux2_1
X_11975_ clknet_leaf_75_clk net442 net368 VGND VGND VPWR VPWR u_decod.pc_q_o\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10926_ u_rf.reg21_q\[16\] _04972_ _05308_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10857_ u_rf.reg20_q\[16\] _04972_ _05271_ VGND VGND VPWR VPWR _05278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10788_ _05241_ VGND VGND VPWR VPWR _00623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12527_ clknet_leaf_38_clk _00564_ net274 VGND VGND VPWR VPWR u_rf.reg17_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ clknet_leaf_24_clk _00495_ net266 VGND VGND VPWR VPWR u_rf.reg15_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11409_ _05570_ VGND VGND VPWR VPWR _00915_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12389_ clknet_leaf_122_clk _00426_ net241 VGND VGND VPWR VPWR u_rf.reg13_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06950_ _01757_ _02044_ _02145_ _01479_ VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a211o_1
X_05901_ u_decod.pc0_q_i\[30\] _01189_ VGND VGND VPWR VPWR _01193_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06881_ _02084_ _02090_ _01744_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_128_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08620_ _03796_ _03798_ _03800_ _03802_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__or4_1
X_05832_ _01139_ _01106_ _01140_ VGND VGND VPWR VPWR _01141_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_124_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08551_ u_rf.reg16_q\[18\] _03323_ _03328_ u_rf.reg12_q\[18\] _03736_ VGND VGND VPWR
+ VPWR _03737_ sky130_fd_sc_hd__a221o_1
X_05763_ u_decod.dec0.instr_i\[4\] _01074_ VGND VGND VPWR VPWR _01086_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_38_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_141_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08482_ u_rf.reg22_q\[15\] _03409_ _03410_ u_rf.reg3_q\[15\] VGND VGND VPWR VPWR
+ _03671_ sky130_fd_sc_hd__a22o_1
X_07502_ _01425_ _02728_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__nand2_1
X_07433_ u_rf.reg0_q\[20\] _01663_ _02371_ u_rf.reg15_q\[20\] _02662_ VGND VGND VPWR
+ VPWR _02663_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09103_ u_decod.pc_q_o\[7\] u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _04238_
+ sky130_fd_sc_hd__nor2_1
X_07364_ u_rf.reg30_q\[19\] _01580_ _01636_ u_rf.reg9_q\[19\] _02595_ VGND VGND VPWR
+ VPWR _02596_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07295_ _02486_ _02488_ _01744_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06315_ _01513_ _01515_ _01566_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__and3_2
XFILLER_0_143_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09034_ _01340_ _01330_ _01337_ _01419_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__or4b_2
X_06246_ _01513_ _01514_ _01515_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__and3_4
XFILLER_0_5_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06177_ u_decod.rs1_data_q\[3\] u_decod.rs1_data_q\[11\] _01376_ u_decod.rs1_data_q\[27\]
+ _01444_ _01447_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09936_ _04767_ VGND VGND VPWR VPWR _00245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09867_ _04422_ _04568_ _04645_ VGND VGND VPWR VPWR _04720_ sky130_fd_sc_hd__or3b_1
X_08818_ u_rf.reg1_q\[30\] _03231_ _03232_ u_rf.reg14_q\[30\] VGND VGND VPWR VPWR
+ _03992_ sky130_fd_sc_hd__a22o_1
X_09798_ _04643_ _04682_ _04645_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__and3_4
X_08749_ u_rf.reg15_q\[27\] _03373_ _03374_ u_rf.reg24_q\[27\] _03925_ VGND VGND VPWR
+ VPWR _03926_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11760_ clknet_leaf_37_clk _00052_ net272 VGND VGND VPWR VPWR u_rf.reg1_q\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ u_rf.reg18_q\[11\] _04962_ _05199_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__mux2_1
X_11691_ _05720_ VGND VGND VPWR VPWR _01047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10642_ _05164_ VGND VGND VPWR VPWR _00554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ u_rf.reg16_q\[10\] _04959_ _05127_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12312_ clknet_leaf_53_clk _00349_ net304 VGND VGND VPWR VPWR u_rf.reg10_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
Xrebuffer9 _04077_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12243_ clknet_leaf_51_clk _00280_ net304 VGND VGND VPWR VPWR u_rf.reg8_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ clknet_leaf_29_clk _00211_ net256 VGND VGND VPWR VPWR u_rf.reg6_q\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11125_ _05420_ VGND VGND VPWR VPWR _00781_ sky130_fd_sc_hd__clkbuf_1
X_11056_ _04749_ u_rf.reg23_q\[13\] _05380_ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__mux2_1
X_10007_ u_rf.reg8_q\[18\] _04465_ _04801_ VGND VGND VPWR VPWR _04810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11958_ clknet_leaf_101_clk net475 net338 VGND VGND VPWR VPWR u_decod.pc_q_o\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11889_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[10\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[10\] sky130_fd_sc_hd__dfrtp_1
X_10909_ u_rf.reg21_q\[8\] _04955_ _05297_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06100_ u_decod.rs1_data_q\[22\] VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_95_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07080_ u_rf.reg17_q\[13\] _01631_ _01791_ u_rf.reg10_q\[13\] _02323_ VGND VGND VPWR
+ VPWR _02324_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06031_ u_decod.rs1_data_q\[10\] VGND VGND VPWR VPWR _01302_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07982_ u_decod.dec0.instr_i\[19\] VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09721_ _04640_ VGND VGND VPWR VPWR _00157_ sky130_fd_sc_hd__clkbuf_1
X_06933_ _01300_ _01429_ _01435_ _01342_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_143_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09652_ _04603_ VGND VGND VPWR VPWR _00125_ sky130_fd_sc_hd__clkbuf_1
X_06864_ u_rf.reg14_q\[9\] _01657_ _01669_ u_rf.reg27_q\[9\] VGND VGND VPWR VPWR _02116_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08603_ u_rf.reg16_q\[20\] _03450_ _03515_ u_rf.reg5_q\[20\] VGND VGND VPWR VPWR
+ _03787_ sky130_fd_sc_hd__a22o_1
X_09583_ u_rf.reg0_q\[30\] _04490_ _04532_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__mux2_1
X_05815_ u_decod.pc0_q_i\[9\] net392 _01127_ VGND VGND VPWR VPWR _01128_ sky130_fd_sc_hd__a21oi_1
X_06795_ u_decod.unsign_ext_q_o net62 net98 VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__and3b_1
X_08534_ u_rf.reg7_q\[17\] _03314_ _03315_ u_rf.reg25_q\[17\] _03720_ VGND VGND VPWR
+ VPWR _03721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05746_ _01068_ _01069_ VGND VGND VPWR VPWR _01070_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08465_ u_rf.reg8_q\[14\] _03270_ _03272_ u_rf.reg29_q\[14\] _03654_ VGND VGND VPWR
+ VPWR _03655_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07416_ _02645_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08396_ u_rf.reg4_q\[11\] _03356_ _03357_ u_rf.reg17_q\[11\] VGND VGND VPWR VPWR
+ _03589_ sky130_fd_sc_hd__a22o_1
X_07347_ _02405_ _02579_ _01472_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_154_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09017_ _04161_ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__nand2_1
X_07278_ u_rf.reg7_q\[17\] _01560_ _01641_ u_rf.reg26_q\[17\] VGND VGND VPWR VPWR
+ _02514_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06229_ _01450_ _01496_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__nand2_4
XFILLER_0_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold150 u_rf.reg12_q\[17\] VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_57_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09919_ _04755_ u_rf.reg7_q\[16\] _04743_ VGND VGND VPWR VPWR _04756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ clknet_leaf_129_clk _00967_ net234 VGND VGND VPWR VPWR u_rf.reg30_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12861_ clknet_leaf_16_clk _00898_ net250 VGND VGND VPWR VPWR u_rf.reg28_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_11812_ clknet_leaf_112_clk net30 net321 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12792_ clknet_leaf_67_clk _00829_ net349 VGND VGND VPWR VPWR u_rf.reg25_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11743_ clknet_leaf_123_clk _00035_ net243 VGND VGND VPWR VPWR u_rf.reg1_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11674_ _05700_ _02418_ _05711_ VGND VGND VPWR VPWR _01039_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10625_ _05155_ VGND VGND VPWR VPWR _00546_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10556_ u_rf.reg16_q\[2\] _04943_ _05116_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10487_ _05081_ VGND VGND VPWR VPWR _00482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12226_ clknet_leaf_130_clk _00263_ net229 VGND VGND VPWR VPWR u_rf.reg8_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12157_ clknet_leaf_14_clk _00194_ net244 VGND VGND VPWR VPWR u_rf.reg6_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_11108_ _05411_ VGND VGND VPWR VPWR _00773_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12088_ clknet_leaf_57_clk _00125_ net292 VGND VGND VPWR VPWR u_rf.reg3_q\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11039_ _04732_ u_rf.reg23_q\[5\] _05369_ VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06580_ u_rf.reg31_q\[3\] _01615_ _01673_ u_rf.reg2_q\[3\] VGND VGND VPWR VPWR _01844_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08250_ _03322_ VGND VGND VPWR VPWR _03450_ sky130_fd_sc_hd__buf_6
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07201_ _02394_ _02396_ _01744_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__o21a_1
X_08181_ u_rf.reg28_q\[2\] _03331_ _03333_ u_rf.reg2_q\[2\] VGND VGND VPWR VPWR _03383_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07132_ _02362_ _02366_ _02370_ _02373_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__or4_1
XFILLER_0_6_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07063_ _01565_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__buf_6
XFILLER_0_140_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06014_ u_decod.rs2_data_q\[26\] u_decod.rs1_data_q\[26\] VGND VGND VPWR VPWR _01285_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07965_ _03170_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__buf_2
X_09704_ u_rf.reg4_q\[21\] _04472_ _04630_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06916_ u_rf.reg31_q\[10\] _01614_ _01648_ u_rf.reg4_q\[10\] VGND VGND VPWR VPWR
+ _02166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ u_rf.reg3_q\[21\] _04472_ _04593_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__mux2_1
X_07896_ u_rf.reg18_q\[30\] _01787_ _02368_ u_rf.reg26_q\[30\] VGND VGND VPWR VPWR
+ _03106_ sky130_fd_sc_hd__a22o_1
X_06847_ _02098_ _02099_ _01444_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__mux2_1
X_09566_ _04557_ VGND VGND VPWR VPWR _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06778_ u_decod.dec0.funct7\[2\] _01530_ _01549_ u_decod.rf_ff_res_data_i\[7\] _02033_
+ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_43_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09497_ _04520_ VGND VGND VPWR VPWR _00053_ sky130_fd_sc_hd__clkbuf_1
X_05729_ u_exe.flush_v_dly1_q u_decod.flush_v VGND VGND VPWR VPWR _01056_ sky130_fd_sc_hd__nor2_4
X_08517_ u_rf.reg27_q\[16\] _03319_ _03321_ u_rf.reg19_q\[16\] _03704_ VGND VGND VPWR
+ VPWR _03705_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_156_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08448_ u_rf.reg3_q\[13\] _03276_ _03556_ u_rf.reg28_q\[13\] _03638_ VGND VGND VPWR
+ VPWR _03639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_147_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10410_ _04786_ u_rf.reg13_q\[31\] _05005_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08379_ u_rf.reg9_q\[10\] _03294_ _03296_ u_rf.reg20_q\[10\] _03572_ VGND VGND VPWR
+ VPWR _03573_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11390_ u_rf.reg28_q\[10\] net505 _05560_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__mux2_1
X_10341_ u_decod.rf_ff_res_data_i\[31\] VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__buf_2
XFILLER_0_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_52_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10272_ _04956_ VGND VGND VPWR VPWR _00392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12011_ clknet_leaf_76_clk u_exe.bu_pc_res\[24\] net369 VGND VGND VPWR VPWR u_exe.pc_data_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ clknet_leaf_22_clk _00950_ net285 VGND VGND VPWR VPWR u_rf.reg29_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_103_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ clknet_leaf_10_clk _00881_ net225 VGND VGND VPWR VPWR u_rf.reg27_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12775_ clknet_leaf_4_clk _00812_ net211 VGND VGND VPWR VPWR u_rf.reg25_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11726_ clknet_leaf_6_clk _00018_ net215 VGND VGND VPWR VPWR u_rf.reg2_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11657_ _05693_ u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10608_ u_rf.reg16_q\[27\] _04995_ _05138_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11588_ _05665_ VGND VGND VPWR VPWR _00999_ sky130_fd_sc_hd__clkbuf_1
X_10539_ _05108_ VGND VGND VPWR VPWR _00507_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_675 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12209_ clknet_leaf_53_clk _00246_ net302 VGND VGND VPWR VPWR u_rf.reg7_q\[22\] sky130_fd_sc_hd__dfrtp_1
X_07750_ u_decod.rs2_data_q\[27\] u_decod.rs1_data_q\[27\] _02781_ VGND VGND VPWR
+ VPWR _02967_ sky130_fd_sc_hd__and3_1
X_06701_ net61 _01487_ _01488_ net47 _01959_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__a221o_1
X_07681_ u_rf.reg11_q\[25\] _01584_ _01595_ u_rf.reg19_q\[25\] _02900_ VGND VGND VPWR
+ VPWR _02901_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09420_ u_rf.reg2_q\[22\] _04474_ _04470_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__mux2_1
X_06632_ u_decod.rf_ff_res_data_i\[4\] _01549_ _01714_ _01874_ _01893_ VGND VGND VPWR
+ VPWR _01894_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09351_ _04427_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__buf_6
XFILLER_0_59_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06563_ net58 _01487_ _01488_ net43 _01827_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08302_ u_decod.pc0_q_i\[6\] _03259_ _03499_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[6\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_23_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ _04385_ _01466_ _04386_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_138_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06494_ net34 _01489_ _01490_ net51 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08233_ u_decod.exe_ff_res_data_i\[3\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[3\]
+ _03433_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08164_ u_rf.reg16_q\[1\] _03322_ _03324_ u_rf.reg5_q\[1\] VGND VGND VPWR VPWR _03367_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_151_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07115_ _01772_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__buf_2
X_08095_ _03269_ _03279_ _03288_ _03298_ VGND VGND VPWR VPWR _03299_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07046_ _02240_ _02290_ _01422_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_149_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08997_ _04144_ _04145_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__xor2_1
X_07948_ u_rf.reg1_q\[31\] _02604_ _02367_ u_rf.reg14_q\[31\] _03155_ VGND VGND VPWR
+ VPWR _03156_ sky130_fd_sc_hd__a221o_1
X_07879_ u_decod.rs1_data_q\[30\] _01371_ _01292_ u_decod.rs1_data_q\[6\] _01469_
+ _01466_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__mux4_1
X_09618_ u_rf.reg3_q\[13\] _04455_ _04582_ VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__mux2_1
X_10890_ u_decod.rf_ff_rd_adr_q_i\[4\] u_decod.rf_write_v_q_i VGND VGND VPWR VPWR
+ _05295_ sky130_fd_sc_hd__and2_1
X_09549_ _04548_ VGND VGND VPWR VPWR _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12560_ clknet_leaf_34_clk _00597_ net269 VGND VGND VPWR VPWR u_rf.reg18_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11511_ _04728_ u_rf.reg30_q\[3\] _05621_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__mux2_1
X_12491_ clknet_leaf_0_clk _00528_ net208 VGND VGND VPWR VPWR u_rf.reg16_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11442_ _05588_ VGND VGND VPWR VPWR _00930_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11373_ u_rf.reg28_q\[2\] net504 _05549_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10324_ u_rf.reg12_q\[25\] _04991_ _04981_ VGND VGND VPWR VPWR _04992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10255_ u_decod.rf_ff_res_data_i\[3\] VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__buf_2
X_10186_ _04732_ u_rf.reg11_q\[5\] _04900_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__mux2_1
Xfanout290 net310 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_85_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12827_ clknet_leaf_10_clk _00864_ net224 VGND VGND VPWR VPWR u_rf.reg27_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12758_ clknet_leaf_48_clk _00795_ net307 VGND VGND VPWR VPWR u_rf.reg24_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12689_ clknet_leaf_55_clk _00726_ net296 VGND VGND VPWR VPWR u_rf.reg22_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11709_ clknet_leaf_108_clk _00001_ net236 VGND VGND VPWR VPWR u_rf.reg2_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08920_ _01289_ u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08851_ _04014_ _04016_ _04013_ VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_0_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07802_ net133 _03007_ _03016_ VGND VGND VPWR VPWR _03017_ sky130_fd_sc_hd__a21o_1
X_08782_ u_rf.reg23_q\[29\] _03354_ _03311_ u_rf.reg1_q\[29\] _03956_ VGND VGND VPWR
+ VPWR _03957_ sky130_fd_sc_hd__a221o_1
X_05994_ u_decod.rs2_data_q\[28\] u_decod.rs1_data_q\[28\] VGND VGND VPWR VPWR _01265_
+ sky130_fd_sc_hd__nor2_1
X_07733_ u_decod.rf_ff_res_data_i\[26\] _02358_ _02743_ _02930_ _02950_ VGND VGND
+ VPWR VPWR _02951_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_79_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07664_ u_decod.dec0.funct7\[0\] _01206_ _02646_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09403_ u_decod.rf_ff_res_data_i\[17\] VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06615_ u_rf.reg30_q\[4\] _01579_ _01624_ u_rf.reg28_q\[4\] VGND VGND VPWR VPWR _01877_
+ sky130_fd_sc_hd__a22o_1
X_07595_ _01368_ _02817_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_9_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09334_ _04409_ u_decod.rs2_data_q\[28\] _04410_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06546_ _01313_ _01319_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__nor2_1
X_09265_ u_decod.pc_q_o\[30\] u_decod.branch_imm_q_o\[30\] VGND VGND VPWR VPWR _04377_
+ sky130_fd_sc_hd__or2_1
X_06477_ u_decod.rs2_data_nxt\[0\] _01744_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__nand2_1
X_09196_ u_decod.pc_q_o\[20\] u_decod.branch_imm_q_o\[20\] VGND VGND VPWR VPWR _04318_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08216_ u_rf.reg26_q\[3\] _03344_ _03345_ u_rf.reg21_q\[3\] VGND VGND VPWR VPWR _03417_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08147_ u_rf.reg9_q\[1\] _03348_ _03349_ u_rf.reg20_q\[1\] VGND VGND VPWR VPWR _03350_
+ sky130_fd_sc_hd__a22o_1
X_08078_ _03202_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__buf_8
XFILLER_0_3_580 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07029_ _02268_ _02270_ _02272_ _02274_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10040_ _04828_ VGND VGND VPWR VPWR _00288_ sky130_fd_sc_hd__clkbuf_1
Xhold65 u_decod.pc0_q_i\[23\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 u_decod.pc0_q_i\[17\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 u_decod.pc0_q_i\[13\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__buf_1
XFILLER_0_98_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11991_ clknet_leaf_87_clk u_exe.bu_pc_res\[4\] net361 VGND VGND VPWR VPWR u_exe.pc_data_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold98 u_decod.pc0_q_i\[5\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlygate4sd3_1
X_10942_ _05323_ VGND VGND VPWR VPWR _00695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10873_ _05286_ VGND VGND VPWR VPWR _00663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ clknet_leaf_110_clk _00649_ net316 VGND VGND VPWR VPWR u_rf.reg20_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12543_ clknet_leaf_132_clk _00580_ net228 VGND VGND VPWR VPWR u_rf.reg18_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12474_ clknet_leaf_94_clk _00511_ net339 VGND VGND VPWR VPWR u_rf.reg15_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11425_ u_rf.reg28_q\[27\] u_decod.rf_ff_res_data_i\[27\] _05571_ VGND VGND VPWR
+ VPWR _05579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 _01579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11356_ _05542_ VGND VGND VPWR VPWR _00890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10307_ u_decod.rf_ff_res_data_i\[20\] VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__buf_2
X_11287_ u_rf.reg26_q\[26\] u_decod.rf_ff_res_data_i\[26\] _05499_ VGND VGND VPWR
+ VPWR _05506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _04784_ u_rf.reg11_q\[30\] _04899_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__mux2_1
X_10169_ u_rf.reg10_q\[30\] _04490_ _04862_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer19 _01060_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_1
XFILLER_0_16_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06400_ _01669_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__buf_6
XFILLER_0_9_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07380_ u_rf.reg19_q\[19\] _01595_ _01791_ u_rf.reg10_q\[19\] _02611_ VGND VGND VPWR
+ VPWR _02612_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_512 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06331_ _01600_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_33_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06262_ u_decod.rf_ff_rd_adr_q_i\[2\] VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__inv_2
X_09050_ _01430_ _04176_ _04191_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08001_ u_rf.reg26_q\[31\] _03203_ _03206_ u_rf.reg21_q\[31\] VGND VGND VPWR VPWR
+ _03207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06193_ _01451_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09952_ u_decod.rf_ff_res_data_i\[27\] VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08903_ _04062_ _04065_ VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09883_ _04731_ VGND VGND VPWR VPWR _00228_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_146_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ u_decod.rs1_data_q\[3\] u_decod.branch_imm_q_o\[3\] VGND VGND VPWR VPWR _04006_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08765_ u_rf.reg31_q\[28\] _03504_ _03505_ u_rf.reg11_q\[28\] _03940_ VGND VGND VPWR
+ VPWR _03941_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07716_ u_rf.reg10_q\[26\] _02380_ _02386_ u_rf.reg27_q\[26\] _02933_ VGND VGND VPWR
+ VPWR _02934_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05977_ _01080_ u_decod.dec0.instr_i\[4\] VGND VGND VPWR VPWR _01252_ sky130_fd_sc_hd__nor2_1
X_08696_ net442 _03773_ _03875_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[24\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07647_ u_decod.pc_q_o\[24\] u_decod.pc_q_o\[25\] _02773_ VGND VGND VPWR VPWR _02868_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_94_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07578_ u_rf.reg16_q\[23\] _01565_ _01631_ u_rf.reg17_q\[23\] VGND VGND VPWR VPWR
+ _02802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09317_ _04406_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
X_06529_ u_rf.reg11_q\[2\] _01584_ _01667_ u_rf.reg8_q\[2\] _01794_ VGND VGND VPWR
+ VPWR _01795_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_62_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09248_ _04328_ _04331_ _04336_ _04361_ _04335_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__a311o_1
XFILLER_0_91_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09179_ _04296_ _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11210_ _05465_ VGND VGND VPWR VPWR _00821_ sky130_fd_sc_hd__clkbuf_1
X_12190_ clknet_leaf_134_clk _00227_ net232 VGND VGND VPWR VPWR u_rf.reg7_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_11141_ u_rf.reg24_q\[21\] _04983_ _05427_ VGND VGND VPWR VPWR _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11072_ _05392_ VGND VGND VPWR VPWR _00756_ sky130_fd_sc_hd__clkbuf_1
Xoutput99 net99 VGND VGND VPWR VPWR access_size_o[1] sky130_fd_sc_hd__buf_2
X_10023_ _04818_ VGND VGND VPWR VPWR _00281_ sky130_fd_sc_hd__clkbuf_1
X_11974_ clknet_leaf_80_clk net439 net371 VGND VGND VPWR VPWR u_decod.pc_q_o\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10925_ _05314_ VGND VGND VPWR VPWR _00687_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10856_ _05277_ VGND VGND VPWR VPWR _00655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_609 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10787_ u_rf.reg19_q\[15\] _04970_ _05235_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12526_ clknet_leaf_28_clk _00563_ net256 VGND VGND VPWR VPWR u_rf.reg17_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ clknet_leaf_21_clk _00494_ net286 VGND VGND VPWR VPWR u_rf.reg15_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_97_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11408_ u_rf.reg28_q\[19\] u_decod.rf_ff_res_data_i\[19\] _05560_ VGND VGND VPWR
+ VPWR _05570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_615 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12388_ clknet_leaf_112_clk _00425_ net317 VGND VGND VPWR VPWR u_rf.reg13_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11339_ _05533_ VGND VGND VPWR VPWR _00882_ sky130_fd_sc_hd__clkbuf_1
X_13009_ clknet_leaf_65_clk _01046_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[22\]
+ sky130_fd_sc_hd__dfxtp_1
X_05900_ u_decod.pc0_q_i\[29\] u_decod.pc0_q_i\[30\] _01186_ VGND VGND VPWR VPWR _01192_
+ sky130_fd_sc_hd__and3_1
X_06880_ _01713_ u_decod.exe_ff_res_data_i\[9\] _02131_ VGND VGND VPWR VPWR _02132_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_128_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05831_ u_decod.pc0_q_i\[11\] u_decod.pc0_q_i\[12\] net411 u_decod.pc0_q_i\[13\]
+ VGND VGND VPWR VPWR _01140_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08550_ u_rf.reg27_q\[18\] _03246_ _03289_ u_rf.reg31_q\[18\] VGND VGND VPWR VPWR
+ _03736_ sky130_fd_sc_hd__a22o_1
X_05762_ _01076_ _01077_ VGND VGND VPWR VPWR _01085_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_141_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08481_ _03197_ VGND VGND VPWR VPWR _03670_ sky130_fd_sc_hd__clkbuf_4
X_07501_ _02724_ _02727_ _02681_ VGND VGND VPWR VPWR _02728_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07432_ u_rf.reg7_q\[20\] _01561_ _01606_ u_rf.reg3_q\[20\] VGND VGND VPWR VPWR _02662_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_99_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09102_ _04029_ _04207_ _04208_ _04237_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[6\]
+ sky130_fd_sc_hd__a2bb2o_1
X_07363_ u_rf.reg2_q\[19\] _01673_ _01666_ u_rf.reg8_q\[19\] VGND VGND VPWR VPWR _02595_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07294_ _01772_ u_decod.exe_ff_res_data_i\[17\] _02529_ VGND VGND VPWR VPWR _02530_
+ sky130_fd_sc_hd__a21o_1
X_06314_ _01583_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09033_ _01420_ _01421_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__and2_1
X_06245_ u_decod.dec0.instr_i\[22\] u_decod.dec0.instr_i\[23\] VGND VGND VPWR VPWR
+ _01515_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06176_ _01446_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09935_ _04766_ u_rf.reg7_q\[21\] _04764_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__mux2_1
X_09866_ u_decod.rf_ff_res_data_i\[0\] VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__buf_2
X_08817_ u_rf.reg15_q\[30\] _03300_ _03302_ u_rf.reg24_q\[30\] _03990_ VGND VGND VPWR
+ VPWR _03991_ sky130_fd_sc_hd__a221o_1
X_09797_ u_decod.rf_ff_rd_adr_q_i\[0\] _01542_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__nor2_1
X_08748_ u_rf.reg6_q\[27\] _03304_ _03306_ u_rf.reg13_q\[27\] VGND VGND VPWR VPWR
+ _03925_ sky130_fd_sc_hd__a22o_1
X_08679_ u_rf.reg8_q\[24\] _03271_ _03273_ u_rf.reg29_q\[24\] _03858_ VGND VGND VPWR
+ VPWR _03859_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_862 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10710_ _05200_ VGND VGND VPWR VPWR _00586_ sky130_fd_sc_hd__clkbuf_1
X_11690_ u_decod.branch_imm_q_o\[23\] _02792_ _05717_ VGND VGND VPWR VPWR _05720_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10641_ u_rf.reg17_q\[10\] _04959_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10572_ _05115_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__buf_6
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12311_ clknet_leaf_71_clk _00348_ net353 VGND VGND VPWR VPWR u_rf.reg10_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12242_ clknet_leaf_40_clk _00279_ net278 VGND VGND VPWR VPWR u_rf.reg8_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12173_ clknet_leaf_6_clk _00210_ net216 VGND VGND VPWR VPWR u_rf.reg6_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11124_ u_rf.reg24_q\[13\] _04966_ _05416_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__mux2_1
X_11055_ _05383_ VGND VGND VPWR VPWR _00748_ sky130_fd_sc_hd__clkbuf_1
X_10006_ _04809_ VGND VGND VPWR VPWR _00273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ clknet_leaf_101_clk net497 net338 VGND VGND VPWR VPWR u_decod.pc_q_o\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_35_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10908_ _05305_ VGND VGND VPWR VPWR _00679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11888_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[9\] net334 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10839_ _05268_ VGND VGND VPWR VPWR _00647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12509_ clknet_leaf_10_clk _00546_ net224 VGND VGND VPWR VPWR u_rf.reg17_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06030_ u_decod.rs2_data_q\[11\] u_decod.rs1_data_q\[11\] VGND VGND VPWR VPWR _01301_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07981_ _03186_ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__inv_2
X_09720_ u_rf.reg4_q\[29\] _04488_ _04630_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__mux2_1
X_06932_ _02180_ _01342_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_143_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ u_rf.reg3_q\[29\] _04488_ _04593_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__mux2_1
X_06863_ u_rf.reg25_q\[9\] _01574_ _01620_ u_rf.reg24_q\[9\] _02114_ VGND VGND VPWR
+ VPWR _02115_ sky130_fd_sc_hd__a221o_1
X_08602_ u_rf.reg7_q\[20\] _03428_ _03429_ u_rf.reg25_q\[20\] _03785_ VGND VGND VPWR
+ VPWR _03786_ sky130_fd_sc_hd__a221o_1
X_09582_ _04565_ VGND VGND VPWR VPWR _00093_ sky130_fd_sc_hd__clkbuf_1
X_05814_ u_decod.pc0_q_i\[9\] net384 _01106_ VGND VGND VPWR VPWR _01127_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06794_ _02048_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__buf_2
X_08533_ u_rf.reg1_q\[17\] _03231_ _03232_ u_rf.reg14_q\[17\] VGND VGND VPWR VPWR
+ _03720_ sky130_fd_sc_hd__a22o_1
X_05745_ u_decod.dec0.instr_i\[0\] u_decod.dec0.instr_i\[1\] u_decod.dec0.instr_i\[2\]
+ VGND VGND VPWR VPWR _01069_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_46_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08464_ u_rf.reg22_q\[14\] _03274_ _03276_ u_rf.reg3_q\[14\] VGND VGND VPWR VPWR
+ _03654_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07415_ u_decod.dec0.funct7\[6\] _02644_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08395_ u_rf.reg8_q\[11\] _03407_ _03408_ u_rf.reg29_q\[11\] _03587_ VGND VGND VPWR
+ VPWR _03588_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07346_ _01468_ _02191_ _01498_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09016_ u_decod.rs1_data_q\[29\] u_decod.branch_imm_q_o\[29\] VGND VGND VPWR VPWR
+ _04162_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07277_ u_rf.reg15_q\[17\] _01600_ _01608_ u_rf.reg12_q\[17\] _02512_ VGND VGND VPWR
+ VPWR _02513_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06228_ _01460_ _01495_ _01498_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold140 u_exe.pc_data_q\[16\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 u_rf.reg28_q\[14\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__dlygate4sd3_1
X_06159_ u_decod.instr_operation_q\[2\] VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_57_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09918_ u_decod.rf_ff_res_data_i\[16\] VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__buf_2
X_09849_ _04710_ VGND VGND VPWR VPWR _00215_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ clknet_leaf_110_clk _00897_ net316 VGND VGND VPWR VPWR u_rf.reg28_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ clknet_leaf_106_clk net29 net319 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_12791_ clknet_leaf_71_clk _00828_ net353 VGND VGND VPWR VPWR u_rf.reg25_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11742_ clknet_leaf_13_clk _00034_ net245 VGND VGND VPWR VPWR u_rf.reg1_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11673_ _05693_ net493 VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10624_ u_rf.reg17_q\[2\] _04943_ _05152_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10555_ _05118_ VGND VGND VPWR VPWR _00513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_40_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10486_ _04726_ u_rf.reg15_q\[2\] _05078_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__mux2_1
X_12225_ clknet_leaf_17_clk _00262_ net251 VGND VGND VPWR VPWR u_rf.reg8_q\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_90_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12156_ clknet_leaf_126_clk _00193_ net239 VGND VGND VPWR VPWR u_rf.reg6_q\[1\] sky130_fd_sc_hd__dfrtp_1
X_11107_ u_rf.reg24_q\[5\] _04949_ _05405_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12087_ clknet_leaf_50_clk _00124_ net308 VGND VGND VPWR VPWR u_rf.reg3_q\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11038_ _05374_ VGND VGND VPWR VPWR _00740_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_121_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12989_ clknet_leaf_92_clk _01026_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08180_ _03197_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__clkbuf_4
X_07200_ _02305_ _02418_ _02439_ VGND VGND VPWR VPWR _02440_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07131_ u_rf.reg15_q\[14\] _02371_ _01610_ u_rf.reg12_q\[14\] _02372_ VGND VGND VPWR
+ VPWR _02373_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07062_ u_decod.dec0.funct3\[1\] _01208_ _02256_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06013_ u_decod.rs2_data_q\[26\] u_decod.rs1_data_q\[26\] VGND VGND VPWR VPWR _01284_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_140_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07964_ u_decod.dec0.instr_i\[19\] VGND VGND VPWR VPWR _03170_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09703_ _04631_ VGND VGND VPWR VPWR _00148_ sky130_fd_sc_hd__clkbuf_1
X_07895_ _01079_ _01224_ _02646_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06915_ _02158_ _02160_ _02162_ _02164_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__or4_1
X_09634_ _04594_ VGND VGND VPWR VPWR _00116_ sky130_fd_sc_hd__clkbuf_1
X_06846_ u_decod.rs1_data_q\[24\] _01702_ _01703_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09565_ u_rf.reg0_q\[21\] _04472_ _04555_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06777_ _01679_ _02032_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__and2_1
X_09496_ u_rf.reg1_q\[21\] _04472_ _04518_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__mux2_1
X_08516_ u_rf.reg16_q\[16\] _03450_ _03515_ u_rf.reg5_q\[16\] VGND VGND VPWR VPWR
+ _03704_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ u_rf.reg7_q\[13\] _03229_ _03230_ u_rf.reg25_q\[13\] VGND VGND VPWR VPWR
+ _03638_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08378_ u_rf.reg31_q\[10\] _03504_ _03505_ u_rf.reg11_q\[10\] VGND VGND VPWR VPWR
+ _03572_ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07329_ u_rf.reg30_q\[18\] _01580_ _01591_ u_rf.reg18_q\[18\] VGND VGND VPWR VPWR
+ _02563_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10340_ _05002_ VGND VGND VPWR VPWR _00414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10271_ u_rf.reg12_q\[8\] _04955_ _04939_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__mux2_1
X_12010_ clknet_leaf_80_clk u_exe.bu_pc_res\[23\] net371 VGND VGND VPWR VPWR u_exe.pc_data_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_72_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12912_ clknet_leaf_36_clk _00949_ net271 VGND VGND VPWR VPWR u_rf.reg29_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_138_clk _00880_ net207 VGND VGND VPWR VPWR u_rf.reg27_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12774_ clknet_leaf_140_clk _00811_ net204 VGND VGND VPWR VPWR u_rf.reg25_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11725_ clknet_leaf_20_clk _00017_ net280 VGND VGND VPWR VPWR u_rf.reg2_q\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_25_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ net457 _05700_ _02644_ _05702_ VGND VGND VPWR VPWR _01030_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10607_ _05145_ VGND VGND VPWR VPWR _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11587_ _04736_ u_rf.reg31_q\[7\] _05657_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10538_ _04778_ u_rf.reg15_q\[27\] _05100_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10469_ _05071_ VGND VGND VPWR VPWR _00474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12208_ clknet_leaf_36_clk _00245_ net273 VGND VGND VPWR VPWR u_rf.reg7_q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12139_ clknet_leaf_0_clk _00176_ net208 VGND VGND VPWR VPWR u_rf.reg5_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_06700_ net38 _01489_ _01490_ net56 VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__a22o_1
X_07680_ u_rf.reg30_q\[25\] _01579_ _01624_ u_rf.reg28_q\[25\] VGND VGND VPWR VPWR
+ _02900_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06631_ _01883_ _01892_ _01679_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__o21a_2
XFILLER_0_87_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09350_ _04423_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__nor2_4
X_06562_ net35 _01489_ _01490_ net52 VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08301_ u_decod.exe_ff_res_data_i\[6\] _03381_ _03498_ VGND VGND VPWR VPWR _03499_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09281_ _04387_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__buf_1
XFILLER_0_142_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06493_ _01480_ _01758_ _01759_ _01442_ VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__o211a_1
X_08232_ _03419_ _03432_ _03337_ VGND VGND VPWR VPWR _03433_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08163_ _03247_ VGND VGND VPWR VPWR _03366_ sky130_fd_sc_hd__buf_8
XFILLER_0_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07114_ _02356_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[14\] sky130_fd_sc_hd__inv_2
XFILLER_0_70_451 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08094_ u_rf.reg31_q\[0\] _03290_ _03292_ u_rf.reg11_q\[0\] _03297_ VGND VGND VPWR
+ VPWR _03298_ sky130_fd_sc_hd__a221o_1
X_07045_ _02193_ _02289_ _01493_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08996_ _04138_ _04140_ _04137_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_149_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07947_ u_rf.reg29_q\[31\] _01780_ _02364_ u_rf.reg21_q\[31\] VGND VGND VPWR VPWR
+ _03155_ sky130_fd_sc_hd__a22o_1
X_07878_ _03052_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09617_ _04585_ VGND VGND VPWR VPWR _00108_ sky130_fd_sc_hd__clkbuf_1
X_06829_ u_decod.dec0.funct7\[3\] _01529_ _01548_ u_decod.rf_ff_res_data_i\[8\] _02082_
+ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09548_ u_rf.reg0_q\[13\] _04455_ _04544_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09479_ u_rf.reg1_q\[13\] _04455_ _04507_ VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11510_ _05624_ VGND VGND VPWR VPWR _00962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12490_ clknet_leaf_29_clk _00527_ net259 VGND VGND VPWR VPWR u_rf.reg16_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11441_ _04726_ u_rf.reg29_q\[2\] _05585_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11372_ _05551_ VGND VGND VPWR VPWR _00897_ sky130_fd_sc_hd__clkbuf_1
X_10323_ u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10254_ _04944_ VGND VGND VPWR VPWR _00386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10185_ _04905_ VGND VGND VPWR VPWR _00356_ sky130_fd_sc_hd__clkbuf_1
Xfanout291 net293 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_4
Xfanout280 net283 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12826_ clknet_leaf_94_clk _00863_ net344 VGND VGND VPWR VPWR u_rf.reg26_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12757_ clknet_leaf_45_clk _00794_ net300 VGND VGND VPWR VPWR u_rf.reg24_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_135_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_135_clk sky130_fd_sc_hd__clkbuf_16
X_12688_ clknet_leaf_32_clk _00725_ net271 VGND VGND VPWR VPWR u_rf.reg22_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11708_ clknet_leaf_11_clk _00000_ net221 VGND VGND VPWR VPWR u_rf.reg2_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11639_ u_decod.dec0.instr_i\[7\] _01227_ _01530_ u_decod.dec0.instr_i\[20\] VGND
+ VGND VPWR VPWR _05692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08850_ _04018_ _04019_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__nor2_1
X_07801_ _01443_ _03011_ _03015_ _01746_ VGND VGND VPWR VPWR _03016_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_71_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08781_ u_rf.reg18_q\[29\] _03222_ _03343_ u_rf.reg26_q\[29\] VGND VGND VPWR VPWR
+ _03956_ sky130_fd_sc_hd__a22o_1
X_05993_ u_decod.rs2_data_q\[28\] u_decod.rs1_data_q\[28\] VGND VGND VPWR VPWR _01264_
+ sky130_fd_sc_hd__and2_1
X_07732_ _02359_ _02949_ VGND VGND VPWR VPWR _02950_ sky130_fd_sc_hd__and2_1
XFILLER_0_149_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07663_ _02332_ _02866_ _02867_ _02883_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[25\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06614_ u_rf.reg25_q\[4\] _01575_ _01622_ u_rf.reg24_q\[4\] _01875_ VGND VGND VPWR
+ VPWR _01876_ sky130_fd_sc_hd__a221o_1
X_09402_ _04462_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__clkbuf_1
X_09333_ _04415_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__dlymetal6s2s_1
X_07594_ _01372_ _01397_ _01369_ _01398_ VGND VGND VPWR VPWR _02817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06545_ _01424_ _01758_ _01809_ _01441_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_126_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_126_clk sky130_fd_sc_hd__clkbuf_16
X_09264_ _04165_ _04206_ _04375_ _04376_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[29\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06476_ _01743_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__inv_2
X_09195_ u_decod.pc_q_o\[20\] u_decod.branch_imm_q_o\[20\] VGND VGND VPWR VPWR _04317_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_118_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08215_ u_rf.reg31_q\[3\] _03290_ _03292_ u_rf.reg11_q\[3\] _03415_ VGND VGND VPWR
+ VPWR _03416_ sky130_fd_sc_hd__a221o_1
X_08146_ _03295_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__buf_8
XFILLER_0_71_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08077_ _03280_ VGND VGND VPWR VPWR _03281_ sky130_fd_sc_hd__buf_8
XFILLER_0_3_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07028_ u_rf.reg20_q\[12\] _01645_ _01671_ u_rf.reg27_q\[12\] _02273_ VGND VGND VPWR
+ VPWR _02274_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08979_ u_decod.rs1_data_q\[24\] u_decod.branch_imm_q_o\[24\] VGND VGND VPWR VPWR
+ _04130_ sky130_fd_sc_hd__nand2_1
Xhold77 u_decod.pc0_q_i\[29\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 u_decod.pc0_q_i\[15\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s25_1
X_11990_ clknet_leaf_89_clk u_exe.bu_pc_res\[3\] net361 VGND VGND VPWR VPWR u_exe.pc_data_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_624 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold99 u_exe.pc_data_q\[8\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 u_decod.exe_ff_rd_adr_q_i\[4\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ u_rf.reg21_q\[23\] _04987_ _05319_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10872_ u_rf.reg20_q\[23\] _04987_ _05282_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_119_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12611_ clknet_leaf_109_clk _00648_ net313 VGND VGND VPWR VPWR u_rf.reg20_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_117_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_117_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12542_ clknet_leaf_134_clk _00579_ net232 VGND VGND VPWR VPWR u_rf.reg18_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12473_ clknet_leaf_57_clk _00510_ net293 VGND VGND VPWR VPWR u_rf.reg15_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11424_ _05578_ VGND VGND VPWR VPWR _00922_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_8 _01581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11355_ _04776_ u_rf.reg27_q\[26\] _05535_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_128_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11286_ _05505_ VGND VGND VPWR VPWR _00857_ sky130_fd_sc_hd__clkbuf_1
X_10306_ _04979_ VGND VGND VPWR VPWR _00403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10237_ _04932_ VGND VGND VPWR VPWR _00381_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10168_ _04895_ VGND VGND VPWR VPWR _00349_ sky130_fd_sc_hd__clkbuf_1
X_10099_ u_rf.reg9_q\[29\] _04488_ _04849_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_137_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_808 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12809_ clknet_leaf_20_clk _00846_ net283 VGND VGND VPWR VPWR u_rf.reg26_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_108_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_108_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06330_ _01599_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06261_ u_decod.rf_ff_rd_adr_q_i\[2\] VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08000_ u_decod.dec0.instr_i\[19\] _03204_ _03205_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__and3_2
XFILLER_0_53_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap200 net201 VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_2
X_06192_ u_decod.rs1_data_q\[6\] _01292_ _01371_ u_decod.rs1_data_q\[30\] _01444_
+ _01447_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09951_ _04777_ VGND VGND VPWR VPWR _00250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08902_ _04050_ _04053_ _04057_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09882_ _04730_ u_rf.reg7_q\[4\] _04722_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ u_decod.rs1_data_q\[3\] u_decod.branch_imm_q_o\[3\] VGND VGND VPWR VPWR _04005_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_146_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ u_rf.reg9_q\[28\] _03293_ _03295_ u_rf.reg20_q\[28\] VGND VGND VPWR VPWR
+ _03940_ sky130_fd_sc_hd__a22o_1
X_05976_ _01251_ VGND VGND VPWR VPWR u_decod.dec0.operation_o\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07715_ u_rf.reg13_q\[26\] _01598_ _02385_ u_rf.reg20_q\[26\] VGND VGND VPWR VPWR
+ _02933_ sky130_fd_sc_hd__a22o_1
X_08695_ u_decod.exe_ff_res_data_i\[24\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[24\]
+ _03874_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07646_ _01277_ _01278_ _02821_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_49_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07577_ _02796_ _02798_ _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__or3_1
XFILLER_0_137_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09316_ _04397_ u_decod.rs2_data_q\[20\] _04398_ VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__and3_1
X_06528_ u_rf.reg1_q\[2\] _01586_ _01636_ u_rf.reg9_q\[2\] VGND VGND VPWR VPWR _01794_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_62_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09247_ _04342_ _04347_ _04360_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_62_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06459_ u_rf.reg24_q\[1\] _01621_ _01627_ u_rf.reg29_q\[1\] VGND VGND VPWR VPWR _01727_
+ sky130_fd_sc_hd__a22o_1
X_09178_ _04283_ _04287_ _04291_ _04297_ _04290_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__a311o_1
X_08129_ _03332_ VGND VGND VPWR VPWR _03333_ sky130_fd_sc_hd__buf_8
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11140_ _05428_ VGND VGND VPWR VPWR _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11071_ _04763_ u_rf.reg23_q\[20\] _05391_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10022_ u_rf.reg8_q\[25\] _04480_ _04812_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__mux2_1
X_11973_ clknet_leaf_80_clk net438 net370 VGND VGND VPWR VPWR u_decod.pc_q_o\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10924_ u_rf.reg21_q\[15\] _04970_ _05308_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10855_ u_rf.reg20_q\[15\] _04970_ _05271_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_587 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10786_ _05240_ VGND VGND VPWR VPWR _00622_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12525_ clknet_leaf_6_clk _00562_ net216 VGND VGND VPWR VPWR u_rf.reg17_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12456_ clknet_leaf_18_clk _00493_ net288 VGND VGND VPWR VPWR u_rf.reg15_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11407_ _05569_ VGND VGND VPWR VPWR _00914_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ clknet_leaf_107_clk _00424_ net315 VGND VGND VPWR VPWR u_rf.reg13_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11338_ _04759_ u_rf.reg27_q\[18\] _05524_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_627 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11269_ _05496_ VGND VGND VPWR VPWR _00849_ sky130_fd_sc_hd__clkbuf_1
X_13008_ clknet_leaf_74_clk _01045_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[21\]
+ sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_145_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05830_ u_decod.pc0_q_i\[12\] u_decod.pc0_q_i\[13\] _01133_ VGND VGND VPWR VPWR _01139_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07500_ _01472_ _02725_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__a21oi_1
X_05761_ _01079_ _01083_ VGND VGND VPWR VPWR _01084_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_141_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ _03187_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_18_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07431_ u_rf.reg29_q\[20\] _01628_ _01639_ u_rf.reg21_q\[20\] _02660_ VGND VGND VPWR
+ VPWR _02661_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07362_ u_decod.dec0.instr_i\[19\] _01208_ _02256_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_459 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09101_ _04233_ _04236_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06313_ _01582_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_154_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07293_ u_decod.rf_ff_res_data_i\[17\] _01549_ _01773_ _02509_ _02528_ VGND VGND
+ VPWR VPWR _02529_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09032_ _04175_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_6
XFILLER_0_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06244_ u_decod.dec0.instr_i\[20\] u_decod.dec0.instr_i\[21\] VGND VGND VPWR VPWR
+ _01514_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06175_ _01445_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09934_ u_decod.rf_ff_res_data_i\[21\] VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09865_ _04718_ VGND VGND VPWR VPWR _00223_ sky130_fd_sc_hd__clkbuf_1
X_08816_ u_rf.reg6_q\[30\] _03235_ _03236_ u_rf.reg13_q\[30\] VGND VGND VPWR VPWR
+ _03990_ sky130_fd_sc_hd__a22o_1
X_09796_ _04681_ VGND VGND VPWR VPWR _00191_ sky130_fd_sc_hd__clkbuf_1
X_08747_ _03917_ _03919_ _03921_ _03923_ VGND VGND VPWR VPWR _03924_ sky130_fd_sc_hd__or4_1
X_05959_ _01238_ VGND VGND VPWR VPWR u_decod.dec0.operation_o\[4\] sky130_fd_sc_hd__clkbuf_1
X_08678_ u_rf.reg22_q\[24\] _03409_ _03277_ u_rf.reg3_q\[24\] VGND VGND VPWR VPWR
+ _03858_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ u_rf.reg21_q\[24\] _01639_ _02386_ u_rf.reg27_q\[24\] VGND VGND VPWR VPWR
+ _02851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10640_ _05151_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__buf_8
XFILLER_0_49_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10571_ _05126_ VGND VGND VPWR VPWR _00521_ sky130_fd_sc_hd__clkbuf_1
X_12310_ clknet_leaf_50_clk _00347_ net308 VGND VGND VPWR VPWR u_rf.reg10_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12241_ clknet_leaf_55_clk _00278_ net294 VGND VGND VPWR VPWR u_rf.reg8_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12172_ clknet_leaf_26_clk _00209_ net266 VGND VGND VPWR VPWR u_rf.reg6_q\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ _05419_ VGND VGND VPWR VPWR _00780_ sky130_fd_sc_hd__clkbuf_1
X_11054_ _04747_ u_rf.reg23_q\[12\] _05380_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__mux2_1
X_10005_ u_rf.reg8_q\[17\] _04463_ _04801_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_106_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11956_ clknet_leaf_100_clk net472 net360 VGND VGND VPWR VPWR u_decod.pc_q_o\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_123_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10907_ u_rf.reg21_q\[7\] _04953_ _05297_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11887_ clknet_leaf_104_clk u_decod.rs2_data_nxt\[8\] net322 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10838_ u_rf.reg20_q\[7\] _04953_ _05260_ VGND VGND VPWR VPWR _05268_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10769_ _05231_ VGND VGND VPWR VPWR _00614_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12508_ clknet_leaf_127_clk _00545_ net237 VGND VGND VPWR VPWR u_rf.reg17_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12439_ clknet_leaf_70_clk _00476_ net353 VGND VGND VPWR VPWR u_rf.reg14_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_752 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07980_ _01257_ _03179_ _03183_ _03185_ VGND VGND VPWR VPWR _03186_ sky130_fd_sc_hd__or4b_1
X_06931_ _01303_ _02134_ VGND VGND VPWR VPWR _02180_ sky130_fd_sc_hd__nand2_1
X_09650_ _04602_ VGND VGND VPWR VPWR _00124_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08601_ u_rf.reg1_q\[20\] _03446_ _03447_ u_rf.reg14_q\[20\] VGND VGND VPWR VPWR
+ _03785_ sky130_fd_sc_hd__a22o_1
X_06862_ u_rf.reg26_q\[9\] _01640_ _01643_ u_rf.reg20_q\[9\] VGND VGND VPWR VPWR _02114_
+ sky130_fd_sc_hd__a22o_1
X_09581_ u_rf.reg0_q\[29\] _04488_ _04555_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__mux2_1
X_05813_ net473 _01105_ _01101_ net95 _01126_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__a221o_1
X_06793_ net99 net112 _01066_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08532_ _03714_ _03716_ _03718_ VGND VGND VPWR VPWR _03719_ sky130_fd_sc_hd__or3_1
X_05744_ u_decod.dec0.instr_i\[4\] u_decod.dec0.instr_i\[5\] u_decod.dec0.instr_i\[6\]
+ VGND VGND VPWR VPWR _01068_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_148_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08463_ u_rf.reg18_q\[14\] _03352_ _03354_ u_rf.reg23_q\[14\] _03652_ VGND VGND VPWR
+ VPWR _03653_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07414_ _02643_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08394_ u_rf.reg22_q\[11\] _03409_ _03410_ u_rf.reg3_q\[11\] VGND VGND VPWR VPWR
+ _03587_ sky130_fd_sc_hd__a22o_1
X_07345_ u_decod.pc_q_o\[18\] u_decod.pc_q_o\[19\] _02506_ VGND VGND VPWR VPWR _02578_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_30_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
X_07276_ u_rf.reg25_q\[17\] _01575_ _01624_ u_rf.reg28_q\[17\] VGND VGND VPWR VPWR
+ _02512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ u_decod.rs1_data_q\[29\] u_decod.branch_imm_q_o\[29\] VGND VGND VPWR VPWR
+ _04161_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06227_ _01497_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold152 u_rf.reg1_q\[23\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 u_exe.pc_data_q\[18\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 u_decod.rf_ff_res_data_i\[2\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__buf_1
X_06158_ _01428_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__buf_4
X_06089_ u_decod.rs2_data_q\[21\] _01358_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_57_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09917_ _04754_ VGND VGND VPWR VPWR _00239_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_97_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
X_09848_ u_rf.reg6_q\[23\] _04476_ _04706_ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ u_rf.reg5_q\[23\] _04476_ _04669_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__mux2_1
X_12790_ clknet_leaf_48_clk _00827_ net306 VGND VGND VPWR VPWR u_rf.reg25_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ clknet_leaf_105_clk net28 net320 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11741_ clknet_leaf_128_clk _00033_ net236 VGND VGND VPWR VPWR u_rf.reg1_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11672_ _05700_ _02391_ _05710_ VGND VGND VPWR VPWR _01038_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10623_ _05154_ VGND VGND VPWR VPWR _00545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_10554_ u_rf.reg16_q\[1\] _04941_ _05116_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10485_ _05080_ VGND VGND VPWR VPWR _00481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12224_ clknet_leaf_119_clk _00261_ net248 VGND VGND VPWR VPWR u_rf.reg8_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12155_ clknet_leaf_10_clk _00192_ net224 VGND VGND VPWR VPWR u_rf.reg6_q\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11106_ _05410_ VGND VGND VPWR VPWR _00772_ sky130_fd_sc_hd__clkbuf_1
X_12086_ clknet_leaf_48_clk _00123_ net306 VGND VGND VPWR VPWR u_rf.reg3_q\[27\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_88_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_125_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11037_ _04730_ u_rf.reg23_q\[4\] _05369_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ clknet_leaf_92_clk _01025_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11939_ clknet_leaf_74_clk u_decod.rs1_data\[27\] net358 VGND VGND VPWR VPWR u_decod.rs1_data_q\[27\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07130_ u_rf.reg25_q\[14\] _01576_ _01625_ u_rf.reg28_q\[14\] VGND VGND VPWR VPWR
+ _02372_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_12_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07061_ _01206_ _01530_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06012_ _01281_ _01282_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_79_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
X_07963_ u_decod.dec0.funct3\[1\] u_decod.dec0.funct3\[2\] _03168_ VGND VGND VPWR
+ VPWR _03169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_156_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09702_ u_rf.reg4_q\[20\] _04469_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__mux2_1
X_07894_ _03104_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[30\] sky130_fd_sc_hd__inv_2
XFILLER_0_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06914_ u_rf.reg5_q\[10\] _01567_ _01594_ u_rf.reg19_q\[10\] _02163_ VGND VGND VPWR
+ VPWR _02164_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09633_ u_rf.reg3_q\[20\] _04469_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__mux2_1
X_06845_ u_decod.rs1_data_q\[16\] _01702_ _01703_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09564_ _04556_ VGND VGND VPWR VPWR _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08515_ u_rf.reg15_q\[16\] _03301_ _03303_ u_rf.reg24_q\[16\] _03702_ VGND VGND VPWR
+ VPWR _03703_ sky130_fd_sc_hd__a221o_1
X_06776_ _02022_ _02031_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09495_ _04519_ VGND VGND VPWR VPWR _00052_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_156_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08446_ u_rf.reg22_q\[13\] _03275_ _03356_ u_rf.reg4_q\[13\] _03636_ VGND VGND VPWR
+ VPWR _03637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08377_ u_rf.reg26_q\[10\] _03344_ _03345_ u_rf.reg21_q\[10\] _03570_ VGND VGND VPWR
+ VPWR _03571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07328_ u_rf.reg17_q\[18\] _01631_ _01791_ u_rf.reg10_q\[18\] _02561_ VGND VGND VPWR
+ VPWR _02562_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07259_ _01757_ _02456_ _02457_ _01423_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10270_ u_decod.rf_ff_res_data_i\[8\] VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_72_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ clknet_leaf_35_clk _00948_ net272 VGND VGND VPWR VPWR u_rf.reg29_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12842_ clknet_leaf_30_clk _00879_ net259 VGND VGND VPWR VPWR u_rf.reg27_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ clknet_leaf_121_clk _00810_ net247 VGND VGND VPWR VPWR u_rf.reg25_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11724_ clknet_leaf_1_clk _00016_ net223 VGND VGND VPWR VPWR u_rf.reg2_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11655_ _05693_ u_decod.branch_imm_q_o\[6\] VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10606_ u_rf.reg16_q\[26\] _04993_ _05138_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__mux2_1
X_11586_ _05664_ VGND VGND VPWR VPWR _00998_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10537_ _05107_ VGND VGND VPWR VPWR _00506_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10468_ _04776_ u_rf.reg14_q\[26\] _05064_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12207_ clknet_leaf_37_clk _00244_ net273 VGND VGND VPWR VPWR u_rf.reg7_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10399_ _05034_ VGND VGND VPWR VPWR _00441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12138_ clknet_leaf_29_clk _00175_ net257 VGND VGND VPWR VPWR u_rf.reg5_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_12069_ clknet_leaf_125_clk _00106_ net239 VGND VGND VPWR VPWR u_rf.reg3_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
X_06630_ _01885_ _01887_ _01889_ _01891_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__or4_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06561_ _01501_ _01706_ _01750_ _01825_ _01479_ _01476_ VGND VGND VPWR VPWR _01826_
+ sky130_fd_sc_hd__mux4_1
X_08300_ u_decod.rf_ff_res_data_i\[6\] _03382_ _03497_ _03404_ VGND VGND VPWR VPWR
+ _03498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06492_ _01424_ _01689_ VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09280_ _04385_ _01469_ _04386_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08231_ _03423_ _03425_ _03427_ _03431_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08162_ _03318_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__buf_8
XFILLER_0_43_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_532 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07113_ _02330_ _02333_ _02337_ _02355_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08093_ u_rf.reg9_q\[0\] _03294_ _03296_ u_rf.reg20_q\[0\] VGND VGND VPWR VPWR _03297_
+ sky130_fd_sc_hd__a22o_1
X_07044_ _02100_ _02288_ _01451_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08995_ _04142_ _04143_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_596 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07946_ u_rf.reg25_q\[31\] _01783_ _01784_ u_rf.reg24_q\[31\] _03153_ VGND VGND VPWR
+ VPWR _03154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07877_ u_decod.instr_operation_q\[0\] u_decod.instr_unit_q\[1\] _01427_ VGND VGND
+ VPWR VPWR _03088_ sky130_fd_sc_hd__nand3_1
XFILLER_0_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06828_ _02072_ _02081_ _01678_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__o21a_1
X_09616_ u_rf.reg3_q\[12\] _04453_ _04582_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__mux2_1
X_09547_ _04547_ VGND VGND VPWR VPWR _00076_ sky130_fd_sc_hd__clkbuf_1
X_06759_ u_rf.reg23_q\[7\] _01612_ _01666_ u_rf.reg8_q\[7\] _02014_ VGND VGND VPWR
+ VPWR _02015_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09478_ _04510_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08429_ u_rf.reg27_q\[12\] _03319_ _03321_ u_rf.reg19_q\[12\] _03620_ VGND VGND VPWR
+ VPWR _03621_ sky130_fd_sc_hd__a221o_1
X_11440_ _05587_ VGND VGND VPWR VPWR _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11371_ u_rf.reg28_q\[1\] net496 _05549_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__mux2_1
X_10322_ _04990_ VGND VGND VPWR VPWR _00408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10253_ u_rf.reg12_q\[2\] _04943_ _04939_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__mux2_1
X_10184_ _04730_ u_rf.reg11_q\[4\] _04900_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__mux2_1
Xfanout292 net293 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout270 net311 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__buf_2
Xfanout281 net283 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12825_ clknet_leaf_64_clk _00862_ net346 VGND VGND VPWR VPWR u_rf.reg26_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12756_ clknet_leaf_30_clk _00793_ net262 VGND VGND VPWR VPWR u_rf.reg24_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12687_ clknet_leaf_42_clk _00724_ net275 VGND VGND VPWR VPWR u_rf.reg22_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11707_ _05728_ VGND VGND VPWR VPWR _01055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11638_ _05691_ VGND VGND VPWR VPWR _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11569_ _04786_ u_rf.reg30_q\[31\] _05620_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08780_ net456 _03773_ _03955_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[28\]
+ sky130_fd_sc_hd__a22o_1
X_07800_ _02965_ _03014_ _01481_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__mux2_1
X_07731_ _02939_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05992_ _01261_ _01262_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07662_ _02868_ _02869_ _02882_ VGND VGND VPWR VPWR _02883_ sky130_fd_sc_hd__o21ai_1
X_07593_ u_decod.pc_q_o\[24\] _02773_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09401_ u_rf.reg2_q\[16\] _04461_ _04449_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__mux2_1
X_06613_ u_rf.reg26_q\[4\] _01641_ _01644_ u_rf.reg20_q\[4\] VGND VGND VPWR VPWR _01875_
+ sky130_fd_sc_hd__a22o_1
X_09332_ _04409_ u_decod.rs2_data_q\[27\] _04410_ VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06544_ _01479_ _01808_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09263_ _04372_ _04373_ _04374_ _04196_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06475_ _01089_ _01739_ _01243_ _01742_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__nor4_2
X_09194_ _04105_ _04274_ _04275_ _04316_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[19\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08214_ u_rf.reg9_q\[3\] _03348_ _03349_ u_rf.reg20_q\[3\] VGND VGND VPWR VPWR _03415_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08145_ _03293_ VGND VGND VPWR VPWR _03348_ sky130_fd_sc_hd__buf_6
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08076_ _03200_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__buf_8
XFILLER_0_101_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07027_ u_rf.reg23_q\[12\] _01612_ _01621_ u_rf.reg24_q\[12\] VGND VGND VPWR VPWR
+ _02273_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08978_ u_decod.rs1_data_q\[24\] u_decod.branch_imm_q_o\[24\] VGND VGND VPWR VPWR
+ _04129_ sky130_fd_sc_hd__or2_1
Xhold78 u_decod.pc0_q_i\[27\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02723_ _03093_ _03137_ _03088_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__a211o_1
Xhold89 _01257_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 u_decod.pc0_q_i\[1\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_2
X_10940_ _05322_ VGND VGND VPWR VPWR _00694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10871_ _05285_ VGND VGND VPWR VPWR _00662_ sky130_fd_sc_hd__clkbuf_1
X_12610_ clknet_leaf_127_clk _00647_ net235 VGND VGND VPWR VPWR u_rf.reg20_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12541_ clknet_leaf_14_clk _00578_ net245 VGND VGND VPWR VPWR u_rf.reg18_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12472_ clknet_leaf_67_clk _00509_ net349 VGND VGND VPWR VPWR u_rf.reg15_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11423_ u_rf.reg28_q\[26\] u_decod.rf_ff_res_data_i\[26\] _05571_ VGND VGND VPWR
+ VPWR _05578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _01581_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11354_ _05541_ VGND VGND VPWR VPWR _00889_ sky130_fd_sc_hd__clkbuf_1
X_11285_ u_rf.reg26_q\[25\] u_decod.rf_ff_res_data_i\[25\] _05499_ VGND VGND VPWR
+ VPWR _05505_ sky130_fd_sc_hd__mux2_1
X_10305_ u_rf.reg12_q\[19\] _04978_ _04960_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10236_ _04782_ u_rf.reg11_q\[29\] _04922_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10167_ u_rf.reg10_q\[29\] _04488_ _04885_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__mux2_1
X_10098_ _04858_ VGND VGND VPWR VPWR _00316_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12808_ clknet_leaf_59_clk _00845_ net290 VGND VGND VPWR VPWR u_rf.reg26_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12739_ clknet_leaf_105_clk _00776_ net320 VGND VGND VPWR VPWR u_rf.reg24_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06260_ _01529_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06191_ u_decod.rs1_data_q\[2\] _01302_ _01384_ u_decod.rs1_data_q\[26\] _01460_
+ _01461_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap201 _01743_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_123_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09950_ _04776_ u_rf.reg7_q\[26\] _04764_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08901_ _01302_ u_decod.branch_imm_q_o\[10\] _04063_ _04056_ VGND VGND VPWR VPWR
+ _04064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09881_ u_decod.rf_ff_res_data_i\[4\] VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__buf_2
XFILLER_0_148_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _03998_ _04004_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_146_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ u_rf.reg18_q\[28\] _03353_ _03355_ u_rf.reg23_q\[28\] _03938_ VGND VGND VPWR
+ VPWR _03939_ sky130_fd_sc_hd__a221o_1
X_05975_ _01227_ _01248_ _01249_ _01250_ VGND VGND VPWR VPWR _01251_ sky130_fd_sc_hd__or4_1
X_07714_ u_rf.reg7_q\[26\] _01562_ _02604_ u_rf.reg1_q\[26\] _02931_ VGND VGND VPWR
+ VPWR _02932_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08694_ _03864_ _03873_ _03378_ VGND VGND VPWR VPWR _03874_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07645_ _01278_ _02821_ _01277_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07576_ u_rf.reg13_q\[23\] _02376_ _01787_ u_rf.reg18_q\[23\] _02799_ VGND VGND VPWR
+ VPWR _02800_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06527_ u_rf.reg23_q\[2\] _01613_ _01791_ u_rf.reg10_q\[2\] _01792_ VGND VGND VPWR
+ VPWR _01793_ sky130_fd_sc_hd__a221o_1
X_09315_ _04405_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_62_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09246_ _04352_ _04355_ _04356_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06458_ _01719_ _01721_ _01723_ _01725_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__or4_1
XFILLER_0_134_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09177_ _04300_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__or2b_1
X_06389_ _01658_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08128_ _03243_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__buf_8
X_08059_ _03223_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__buf_8
X_11070_ _05368_ VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10021_ _04817_ VGND VGND VPWR VPWR _00280_ sky130_fd_sc_hd__clkbuf_1
X_11972_ clknet_leaf_79_clk net443 net370 VGND VGND VPWR VPWR u_decod.pc_q_o\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_488 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10923_ _05313_ VGND VGND VPWR VPWR _00686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10854_ _05276_ VGND VGND VPWR VPWR _00654_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10785_ net523 _04968_ _05235_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12524_ clknet_leaf_9_clk _00561_ net225 VGND VGND VPWR VPWR u_rf.reg17_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_273 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12455_ clknet_leaf_11_clk _00492_ net223 VGND VGND VPWR VPWR u_rf.reg15_q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_113_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11406_ u_rf.reg28_q\[18\] u_decod.rf_ff_res_data_i\[18\] _05560_ VGND VGND VPWR
+ VPWR _05569_ sky130_fd_sc_hd__mux2_1
X_12386_ clknet_leaf_130_clk _00423_ net229 VGND VGND VPWR VPWR u_rf.reg13_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11337_ _05532_ VGND VGND VPWR VPWR _00881_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11268_ u_rf.reg26_q\[17\] u_decod.rf_ff_res_data_i\[17\] _05488_ VGND VGND VPWR
+ VPWR _05496_ sky130_fd_sc_hd__mux2_1
X_10219_ _04923_ VGND VGND VPWR VPWR _00372_ sky130_fd_sc_hd__clkbuf_1
X_13007_ clknet_leaf_65_clk _01044_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[20\]
+ sky130_fd_sc_hd__dfxtp_2
X_11199_ _05459_ VGND VGND VPWR VPWR _00816_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05760_ _01080_ u_decod.dec0.funct7\[6\] _01082_ VGND VGND VPWR VPWR _01083_ sky130_fd_sc_hd__or3_1
XFILLER_0_89_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07430_ u_rf.reg1_q\[20\] _01587_ _01659_ u_rf.reg14_q\[20\] VGND VGND VPWR VPWR
+ _02660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07361_ _02575_ _02576_ _02593_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[19\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09100_ _04223_ _04224_ _04226_ _04234_ _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06312_ _01512_ _01558_ _01573_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__and3_2
XFILLER_0_150_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09031_ net133 _04174_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__and2_4
XFILLER_0_115_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07292_ _02511_ _02520_ _02527_ _01679_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__o31a_2
XFILLER_0_60_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06243_ _01512_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06174_ u_decod.rs2_data_q\[4\] VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09933_ _04765_ VGND VGND VPWR VPWR _00244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09864_ u_rf.reg6_q\[31\] _04492_ _04683_ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08815_ u_rf.reg27_q\[30\] _03318_ _03320_ u_rf.reg19_q\[30\] _03988_ VGND VGND VPWR
+ VPWR _03989_ sky130_fd_sc_hd__a221o_1
X_09795_ u_rf.reg5_q\[31\] _04492_ _04646_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08746_ u_rf.reg30_q\[27\] _03281_ _03283_ u_rf.reg10_q\[27\] _03922_ VGND VGND VPWR
+ VPWR _03923_ sky130_fd_sc_hd__a221o_1
X_05958_ _01205_ _01237_ VGND VGND VPWR VPWR _01238_ sky130_fd_sc_hd__or2_1
X_05889_ u_decod.pc0_q_i\[27\] _01180_ VGND VGND VPWR VPWR _01184_ sky130_fd_sc_hd__nand2_1
X_08677_ u_rf.reg18_q\[24\] _03262_ _03263_ u_rf.reg23_q\[24\] _03856_ VGND VGND VPWR
+ VPWR _03857_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_37_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _02843_ _02845_ _02847_ _02849_ VGND VGND VPWR VPWR _02850_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07559_ _01746_ _02780_ _02783_ _01260_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10570_ u_rf.reg16_q\[9\] _04957_ _05116_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__mux2_1
X_09229_ u_decod.pc_q_o\[25\] u_decod.branch_imm_q_o\[25\] VGND VGND VPWR VPWR _04346_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_91_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12240_ clknet_leaf_34_clk _00277_ net276 VGND VGND VPWR VPWR u_rf.reg8_q\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_79_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12171_ clknet_leaf_0_clk _00208_ net208 VGND VGND VPWR VPWR u_rf.reg6_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11122_ u_rf.reg24_q\[12\] _04964_ _05416_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__mux2_1
X_11053_ _05382_ VGND VGND VPWR VPWR _00747_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10004_ _04808_ VGND VGND VPWR VPWR _00272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11955_ clknet_leaf_86_clk net386 net338 VGND VGND VPWR VPWR u_decod.pc_q_o\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ _05304_ VGND VGND VPWR VPWR _00678_ sky130_fd_sc_hd__clkbuf_1
X_11886_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[7\] net322 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10837_ _05267_ VGND VGND VPWR VPWR _00646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10768_ u_rf.reg19_q\[6\] _04951_ _05224_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12507_ clknet_leaf_12_clk _00544_ net221 VGND VGND VPWR VPWR u_rf.reg17_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_506 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12438_ clknet_leaf_47_clk _00475_ net306 VGND VGND VPWR VPWR u_rf.reg14_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _05194_ VGND VGND VPWR VPWR _00581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12369_ clknet_leaf_56_clk _00406_ net287 VGND VGND VPWR VPWR u_rf.reg12_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06930_ _02177_ _02179_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[10\] sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_143_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ u_rf.reg15_q\[20\] _03373_ _03374_ u_rf.reg24_q\[20\] _03783_ VGND VGND VPWR
+ VPWR _03784_ sky130_fd_sc_hd__a221o_1
X_06861_ u_rf.reg13_q\[9\] _01596_ _01590_ u_rf.reg18_q\[9\] _02112_ VGND VGND VPWR
+ VPWR _02113_ sky130_fd_sc_hd__a221o_1
X_09580_ _04564_ VGND VGND VPWR VPWR _00092_ sky130_fd_sc_hd__clkbuf_1
X_05812_ _01124_ _01106_ _01125_ VGND VGND VPWR VPWR _01126_ sky130_fd_sc_hd__and3b_1
X_06792_ net99 _01064_ _01067_ net100 VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__a31o_2
X_08531_ u_rf.reg8_q\[17\] _03270_ _03272_ u_rf.reg29_q\[17\] _03717_ VGND VGND VPWR
+ VPWR _03718_ sky130_fd_sc_hd__a221o_1
X_05743_ _01067_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__inv_2
XFILLER_0_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08462_ u_rf.reg4_q\[14\] _03264_ _03266_ u_rf.reg17_q\[14\] VGND VGND VPWR VPWR
+ _03652_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07413_ _01226_ _01715_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__or2_1
XFILLER_0_148_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08393_ u_decod.pc0_q_i\[10\] _03565_ _03585_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[10\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07344_ u_decod.pc_q_o\[18\] _02506_ u_decod.pc_q_o\[19\] VGND VGND VPWR VPWR _02577_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07275_ u_rf.reg16_q\[17\] _01565_ _01674_ u_rf.reg2_q\[17\] _02510_ VGND VGND VPWR
+ VPWR _02511_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09014_ _04101_ _04160_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__nor2_1
XFILLER_0_116_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06226_ u_decod.rs2_data_q\[3\] _01496_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__nand2_2
XFILLER_0_103_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold142 u_exe.pc_data_q\[4\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 u_exe.pc_data_q\[1\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 u_decod.rf_ff_res_data_i\[10\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 u_rf.reg24_q\[16\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__dlygate4sd3_1
X_06157_ u_decod.instr_unit_q\[0\] u_decod.instr_operation_q\[1\] _01427_ VGND VGND
+ VPWR VPWR _01428_ sky130_fd_sc_hd__and3_1
X_06088_ u_decod.rs2_data_q\[21\] _01358_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_57_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09916_ _04753_ u_rf.reg7_q\[15\] _04743_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__mux2_1
X_09847_ _04709_ VGND VGND VPWR VPWR _00214_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09778_ _04672_ VGND VGND VPWR VPWR _00182_ sky130_fd_sc_hd__clkbuf_1
X_08729_ u_rf.reg1_q\[26\] _03446_ _03447_ u_rf.reg14_q\[26\] VGND VGND VPWR VPWR
+ _03907_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11740_ clknet_leaf_13_clk _00032_ net245 VGND VGND VPWR VPWR u_rf.reg1_q\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11671_ _05693_ net485 VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10622_ u_rf.reg17_q\[1\] _04941_ _05152_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10553_ _05117_ VGND VGND VPWR VPWR _00512_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10484_ _04724_ u_rf.reg15_q\[1\] _05078_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12223_ clknet_leaf_131_clk _00260_ net227 VGND VGND VPWR VPWR u_rf.reg8_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12154_ clknet_leaf_58_clk _00191_ net292 VGND VGND VPWR VPWR u_rf.reg5_q\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11105_ u_rf.reg24_q\[4\] _04947_ _05405_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__mux2_1
X_12085_ clknet_leaf_47_clk _00122_ net300 VGND VGND VPWR VPWR u_rf.reg3_q\[26\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11036_ _05373_ VGND VGND VPWR VPWR _00739_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12987_ clknet_leaf_92_clk _01024_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[0\]
+ sky130_fd_sc_hd__dfxtp_2
X_11938_ clknet_leaf_74_clk u_decod.rs1_data\[26\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11869_ clknet_leaf_103_clk u_decod.dec0.operation_o\[0\] net335 VGND VGND VPWR VPWR
+ u_decod.instr_operation_q\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_156_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07060_ _01437_ _02282_ _02283_ _02304_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[13\]
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_136_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06011_ u_decod.rs2_data_q\[27\] u_decod.rs1_data_q\[27\] VGND VGND VPWR VPWR _01282_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_70_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09701_ _04607_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__buf_6
X_07962_ _01080_ _01071_ _01075_ _01094_ _01212_ VGND VGND VPWR VPWR _03168_ sky130_fd_sc_hd__a41o_1
XFILLER_0_156_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07893_ _03084_ _03085_ _03103_ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06913_ u_rf.reg16_q\[10\] _01563_ _01629_ u_rf.reg17_q\[10\] VGND VGND VPWR VPWR
+ _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09632_ _04570_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_52_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06844_ _01478_ _02045_ _02096_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__o21ai_1
X_09563_ u_rf.reg0_q\[20\] _04469_ _04555_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08514_ u_rf.reg6_q\[16\] _03305_ _03388_ u_rf.reg13_q\[16\] VGND VGND VPWR VPWR
+ _03702_ sky130_fd_sc_hd__a22o_1
X_06775_ _02024_ _02026_ _02028_ _02030_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__or4_1
X_09494_ net520 _04469_ _04518_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08445_ u_rf.reg10_q\[13\] _03202_ _03332_ u_rf.reg2_q\[13\] VGND VGND VPWR VPWR
+ _03636_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_156_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08376_ u_rf.reg30_q\[10\] _03280_ _03282_ u_rf.reg10_q\[10\] VGND VGND VPWR VPWR
+ _03570_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07327_ u_rf.reg29_q\[18\] _01627_ _01653_ u_rf.reg22_q\[18\] VGND VGND VPWR VPWR
+ _02561_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07258_ _02406_ _02494_ _01757_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07189_ u_rf.reg30_q\[15\] _01580_ _01592_ u_rf.reg18_q\[15\] VGND VGND VPWR VPWR
+ _02429_ sky130_fd_sc_hd__a22o_1
X_06209_ _01479_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ clknet_leaf_28_clk _00947_ net258 VGND VGND VPWR VPWR u_rf.reg29_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12841_ clknet_leaf_22_clk _00878_ net284 VGND VGND VPWR VPWR u_rf.reg27_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_103_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ clknet_leaf_111_clk _00809_ net316 VGND VGND VPWR VPWR u_rf.reg25_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11723_ clknet_leaf_29_clk _00015_ net257 VGND VGND VPWR VPWR u_rf.reg2_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11654_ net458 _05700_ _02644_ _05701_ VGND VGND VPWR VPWR _01029_ sky130_fd_sc_hd__a31o_1
XFILLER_0_154_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10605_ _05144_ VGND VGND VPWR VPWR _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11585_ _04734_ u_rf.reg31_q\[6\] _05657_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10536_ _04776_ u_rf.reg15_q\[26\] _05100_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10467_ _05070_ VGND VGND VPWR VPWR _00473_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12206_ clknet_leaf_27_clk _00243_ net258 VGND VGND VPWR VPWR u_rf.reg7_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10398_ _04774_ u_rf.reg13_q\[25\] _05028_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_575 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12137_ clknet_leaf_24_clk _00174_ net265 VGND VGND VPWR VPWR u_rf.reg5_q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12068_ clknet_leaf_108_clk _00105_ net312 VGND VGND VPWR VPWR u_rf.reg3_q\[9\] sky130_fd_sc_hd__dfrtp_1
X_11019_ u_rf.reg22_q\[28\] _04997_ _05355_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06560_ _01464_ _01824_ _01500_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06491_ _01452_ _01756_ _01757_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08230_ u_rf.reg7_q\[3\] _03428_ _03429_ u_rf.reg25_q\[3\] _03430_ VGND VGND VPWR
+ VPWR _03431_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08161_ u_rf.reg0_q\[1\] _03175_ _03328_ u_rf.reg12_q\[1\] _03363_ VGND VGND VPWR
+ VPWR _03364_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_151_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08092_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__buf_6
X_07112_ _01746_ _02341_ _02354_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_141_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07043_ _02286_ _02287_ _01455_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_599 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08994_ u_decod.rs1_data_q\[26\] u_decod.branch_imm_q_o\[26\] VGND VGND VPWR VPWR
+ _04143_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07945_ u_rf.reg26_q\[31\] _02368_ _02385_ u_rf.reg20_q\[31\] VGND VGND VPWR VPWR
+ _03153_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07876_ u_decod.pc_q_o\[29\] u_decod.pc_q_o\[30\] _02999_ VGND VGND VPWR VPWR _03087_
+ sky130_fd_sc_hd__and3_1
X_09615_ _04584_ VGND VGND VPWR VPWR _00107_ sky130_fd_sc_hd__clkbuf_1
X_06827_ _02074_ _02076_ _02078_ _02080_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__or4_1
X_09546_ u_rf.reg0_q\[12\] _04453_ _04544_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__mux2_1
X_06758_ u_rf.reg11_q\[7\] _01582_ _01634_ u_rf.reg9_q\[7\] VGND VGND VPWR VPWR _02014_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09477_ u_rf.reg1_q\[12\] _04453_ _04507_ VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08428_ u_rf.reg16_q\[12\] _03450_ _03515_ u_rf.reg5_q\[12\] VGND VGND VPWR VPWR
+ _03620_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _01330_ _01947_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08359_ u_rf.reg15_q\[9\] _03300_ _03302_ u_rf.reg24_q\[9\] VGND VGND VPWR VPWR _03554_
+ sky130_fd_sc_hd__a22o_1
X_11370_ _05550_ VGND VGND VPWR VPWR _00896_ sky130_fd_sc_hd__clkbuf_1
X_10321_ u_rf.reg12_q\[24\] _04989_ _04981_ VGND VGND VPWR VPWR _04990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10252_ u_decod.rf_ff_res_data_i\[2\] VGND VGND VPWR VPWR _04943_ sky130_fd_sc_hd__clkbuf_4
X_10183_ _04904_ VGND VGND VPWR VPWR _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout271 net274 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_4
Xfanout282 net283 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout260 net270 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_2
Xfanout293 net310 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_4
X_12824_ clknet_leaf_65_clk _00861_ net355 VGND VGND VPWR VPWR u_rf.reg26_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12755_ clknet_leaf_52_clk _00792_ net304 VGND VGND VPWR VPWR u_rf.reg24_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11706_ u_decod.branch_imm_q_o\[31\] _03143_ net346 VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_658 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12686_ clknet_leaf_28_clk _00723_ net258 VGND VGND VPWR VPWR u_rf.reg22_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11637_ _04786_ u_rf.reg31_q\[31\] _05656_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11568_ _05654_ VGND VGND VPWR VPWR _00990_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10519_ _04759_ u_rf.reg15_q\[18\] _05089_ VGND VGND VPWR VPWR _05098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11499_ _04784_ u_rf.reg29_q\[30\] _05584_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07730_ _02941_ _02943_ _02945_ _02947_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__or4_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05991_ u_decod.rs2_data_q\[29\] u_decod.rs1_data_q\[29\] VGND VGND VPWR VPWR _01262_
+ sky130_fd_sc_hd__and2_1
X_07661_ _02789_ _02873_ _02879_ _02881_ VGND VGND VPWR VPWR _02882_ sky130_fd_sc_hd__o211a_1
X_07592_ u_decod.pc_q_o\[24\] _02773_ VGND VGND VPWR VPWR _02815_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06612_ u_decod.dec0.instr_i\[11\] _01226_ _01715_ _01572_ VGND VGND VPWR VPWR _01874_
+ sky130_fd_sc_hd__a22o_1
X_09400_ u_decod.rf_ff_res_data_i\[16\] VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09331_ _04414_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_1
X_06543_ _01687_ _01807_ _01688_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09262_ _04372_ _04373_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06474_ _01079_ _01075_ _01740_ _01741_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__and4_1
XFILLER_0_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09193_ _04313_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08213_ u_rf.reg18_q\[3\] _03353_ _03355_ u_rf.reg23_q\[3\] _03413_ VGND VGND VPWR
+ VPWR _03414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08144_ u_rf.reg30_q\[1\] _03341_ _03342_ u_rf.reg10_q\[1\] _03346_ VGND VGND VPWR
+ VPWR _03347_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08075_ u_rf.reg8_q\[0\] _03271_ _03273_ u_rf.reg29_q\[0\] _03278_ VGND VGND VPWR
+ VPWR _03279_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07026_ u_rf.reg16_q\[12\] _01565_ _01674_ u_rf.reg2_q\[12\] _02271_ VGND VGND VPWR
+ VPWR _02272_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08977_ _04101_ _04128_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__nor2_1
Xhold68 u_decod.pc0_q_i\[24\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 u_decod.pc0_q_i\[16\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _02723_ _03136_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__nor2_1
X_07859_ u_rf.reg29_q\[29\] _01780_ _01776_ u_rf.reg2_q\[29\] _03070_ VGND VGND VPWR
+ VPWR _03071_ sky130_fd_sc_hd__a221o_1
X_10870_ u_rf.reg20_q\[22\] _04985_ _05282_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09529_ u_rf.reg0_q\[4\] _04436_ _04533_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_320 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12540_ clknet_leaf_127_clk _00577_ net235 VGND VGND VPWR VPWR u_rf.reg18_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12471_ clknet_leaf_70_clk _00508_ net353 VGND VGND VPWR VPWR u_rf.reg15_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11422_ _05577_ VGND VGND VPWR VPWR _00921_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11353_ _04774_ u_rf.reg27_q\[25\] _05535_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11284_ _05504_ VGND VGND VPWR VPWR _00856_ sky130_fd_sc_hd__clkbuf_1
X_10304_ u_decod.rf_ff_res_data_i\[19\] VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__buf_2
X_10235_ _04931_ VGND VGND VPWR VPWR _00380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10166_ _04894_ VGND VGND VPWR VPWR _00348_ sky130_fd_sc_hd__clkbuf_1
X_10097_ u_rf.reg9_q\[28\] _04486_ _04849_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_350 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12807_ clknet_leaf_3_clk _00844_ net213 VGND VGND VPWR VPWR u_rf.reg26_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_10999_ _05353_ VGND VGND VPWR VPWR _00722_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12738_ clknet_leaf_133_clk _00775_ net230 VGND VGND VPWR VPWR u_rf.reg24_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12669_ clknet_leaf_14_clk _00706_ net246 VGND VGND VPWR VPWR u_rf.reg22_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06190_ _01447_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_13_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08900_ u_decod.rs1_data_q\[11\] u_decod.branch_imm_q_o\[11\] VGND VGND VPWR VPWR
+ _04063_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09880_ _04729_ VGND VGND VPWR VPWR _00227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08831_ _04000_ _04003_ VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_146_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ u_rf.reg4_q\[28\] _03265_ _03267_ u_rf.reg17_q\[28\] VGND VGND VPWR VPWR
+ _03938_ sky130_fd_sc_hd__a22o_1
X_05974_ _01075_ _01219_ _01198_ VGND VGND VPWR VPWR _01250_ sky130_fd_sc_hd__and3_1
X_07713_ u_rf.reg15_q\[26\] _01601_ _02363_ u_rf.reg3_q\[26\] VGND VGND VPWR VPWR
+ _02931_ sky130_fd_sc_hd__a22o_1
X_08693_ _03866_ _03868_ _03870_ _03872_ VGND VGND VPWR VPWR _03873_ sky130_fd_sc_hd__or4_1
X_07644_ _02862_ _02865_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[24\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07575_ u_rf.reg23_q\[23\] _02652_ _01791_ u_rf.reg10_q\[23\] VGND VGND VPWR VPWR
+ _02799_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06526_ u_rf.reg6_q\[2\] _01556_ _01653_ u_rf.reg22_q\[2\] VGND VGND VPWR VPWR _01792_
+ sky130_fd_sc_hd__a22o_1
X_09314_ _04397_ u_decod.rs2_data_q\[19\] _04398_ VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and3_1
X_09245_ _04151_ _04206_ _04197_ _04359_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[27\]
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_62_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06457_ u_rf.reg0_q\[1\] _01662_ _01670_ u_rf.reg27_q\[1\] _01724_ VGND VGND VPWR
+ VPWR _01725_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_32_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09176_ u_decod.pc_q_o\[17\] u_decod.branch_imm_q_o\[17\] VGND VGND VPWR VPWR _04301_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06388_ _01657_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__buf_6
XFILLER_0_133_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08127_ _03330_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08058_ _03222_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__buf_8
XFILLER_0_102_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07009_ _02255_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[12\] sky130_fd_sc_hd__buf_1
X_10020_ u_rf.reg8_q\[24\] _04478_ _04812_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__mux2_1
X_11971_ clknet_leaf_80_clk net445 net370 VGND VGND VPWR VPWR u_decod.pc_q_o\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ u_rf.reg21_q\[14\] _04968_ _05308_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10853_ u_rf.reg20_q\[14\] _04968_ _05271_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10784_ _05239_ VGND VGND VPWR VPWR _00621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12523_ clknet_leaf_136_clk _00560_ net205 VGND VGND VPWR VPWR u_rf.reg17_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_285 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12454_ clknet_leaf_138_clk _00491_ net210 VGND VGND VPWR VPWR u_rf.reg15_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11405_ _05568_ VGND VGND VPWR VPWR _00913_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12385_ clknet_leaf_117_clk _00422_ net325 VGND VGND VPWR VPWR u_rf.reg13_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11336_ _04757_ u_rf.reg27_q\[17\] _05524_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13006_ clknet_leaf_65_clk _01043_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[19\]
+ sky130_fd_sc_hd__dfxtp_2
X_11267_ _05495_ VGND VGND VPWR VPWR _00848_ sky130_fd_sc_hd__clkbuf_1
X_10218_ _04763_ u_rf.reg11_q\[20\] _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__mux2_1
X_11198_ u_rf.reg25_q\[16\] _04972_ _05452_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__mux2_1
X_10149_ u_rf.reg10_q\[20\] _04469_ _04885_ VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07360_ _02334_ _02577_ _02578_ _02592_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__o31a_1
XFILLER_0_57_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06311_ _01580_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_44_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09030_ _04172_ _04173_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07291_ _02522_ _02524_ _02526_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06242_ u_decod.dec0.instr_i\[24\] VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06173_ u_decod.rs2_data_q\[3\] VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09932_ _04763_ u_rf.reg7_q\[20\] _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09863_ _04717_ VGND VGND VPWR VPWR _00222_ sky130_fd_sc_hd__clkbuf_1
X_09794_ _04680_ VGND VGND VPWR VPWR _00190_ sky130_fd_sc_hd__clkbuf_1
X_08814_ u_rf.reg16_q\[30\] _03248_ _03249_ u_rf.reg5_q\[30\] VGND VGND VPWR VPWR
+ _03988_ sky130_fd_sc_hd__a22o_1
X_08745_ u_rf.reg26_q\[27\] _03284_ _03286_ u_rf.reg21_q\[27\] VGND VGND VPWR VPWR
+ _03922_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_77_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05957_ _01089_ _01233_ _01236_ VGND VGND VPWR VPWR _01237_ sky130_fd_sc_hd__nand3b_2
X_05888_ u_decod.pc0_q_i\[27\] _01180_ VGND VGND VPWR VPWR _01183_ sky130_fd_sc_hd__or2_1
X_08676_ u_rf.reg4_q\[24\] _03264_ _03266_ u_rf.reg17_q\[24\] VGND VGND VPWR VPWR
+ _03856_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_37_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ u_rf.reg3_q\[24\] _02363_ _02697_ u_rf.reg4_q\[24\] _02848_ VGND VGND VPWR
+ VPWR _02849_ sky130_fd_sc_hd__a221o_1
X_07558_ _02781_ _01369_ _02770_ _01435_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06509_ u_decod.rf_ff_res_data_i\[2\] _01549_ _01773_ _01774_ VGND VGND VPWR VPWR
+ _01775_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07489_ u_decod.rf_ff_res_data_i\[21\] _01550_ _01773_ _02696_ _02716_ VGND VGND
+ VPWR VPWR _02717_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09228_ u_decod.pc_q_o\[25\] u_decod.branch_imm_q_o\[25\] VGND VGND VPWR VPWR _04345_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09159_ _04284_ _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_890 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ clknet_leaf_30_clk _00207_ net261 VGND VGND VPWR VPWR u_rf.reg6_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11121_ _05418_ VGND VGND VPWR VPWR _00779_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11052_ _04745_ u_rf.reg23_q\[11\] _05380_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__mux2_1
X_10003_ u_rf.reg8_q\[16\] _04461_ _04801_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11954_ clknet_leaf_100_clk net389 net338 VGND VGND VPWR VPWR u_decod.pc_q_o\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ u_rf.reg21_q\[6\] _04951_ _05297_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__mux2_1
X_11885_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[6\] net322 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10836_ u_rf.reg20_q\[6\] _04951_ _05260_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10767_ _05230_ VGND VGND VPWR VPWR _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12506_ clknet_leaf_58_clk _00543_ net292 VGND VGND VPWR VPWR u_rf.reg16_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ u_rf.reg18_q\[5\] _04949_ _05188_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12437_ clknet_leaf_47_clk _00474_ net300 VGND VGND VPWR VPWR u_rf.reg14_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12368_ clknet_leaf_35_clk _00405_ net276 VGND VGND VPWR VPWR u_rf.reg12_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11319_ _04740_ u_rf.reg27_q\[9\] _05513_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__mux2_1
X_12299_ clknet_leaf_134_clk _00336_ net209 VGND VGND VPWR VPWR u_rf.reg10_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_06860_ u_rf.reg30_q\[9\] _01578_ _01623_ u_rf.reg28_q\[9\] VGND VGND VPWR VPWR _02112_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05811_ u_decod.pc0_q_i\[8\] _01121_ VGND VGND VPWR VPWR _01125_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06791_ _02002_ _02045_ _01478_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08530_ u_rf.reg22_q\[17\] _03274_ _03276_ u_rf.reg3_q\[17\] VGND VGND VPWR VPWR
+ _03717_ sky130_fd_sc_hd__a22o_1
X_05742_ _01057_ _01066_ VGND VGND VPWR VPWR _01067_ sky130_fd_sc_hd__or2_1
X_08461_ u_rf.reg9_q\[14\] _03348_ _03349_ u_rf.reg20_q\[14\] _03650_ VGND VGND VPWR
+ VPWR _03651_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_46_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07412_ _02642_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[20\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08392_ _03178_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07343_ _01386_ _01379_ _02534_ _01765_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07274_ u_rf.reg1_q\[17\] _01587_ _01667_ u_rf.reg8_q\[17\] VGND VGND VPWR VPWR _02510_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09013_ _04156_ _04159_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06225_ _01267_ _01430_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__nand2_2
Xhold110 u_exe.pc_data_q\[26\] VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 u_exe.pc_data_q\[23\] VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold143 u_exe.pc_data_q\[21\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 u_exe.pc_data_q\[29\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06156_ _01056_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_4
Xhold154 u_rf.reg3_q\[24\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__dlygate4sd3_1
X_06087_ u_decod.rs1_data_q\[21\] VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_57_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09915_ u_decod.rf_ff_res_data_i\[15\] VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__buf_2
X_09846_ u_rf.reg6_q\[22\] _04474_ _04706_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ u_rf.reg5_q\[22\] _04474_ _04669_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__mux2_1
X_06989_ u_decod.rs1_data_q\[19\] _01454_ _01753_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__o21a_1
X_08728_ u_rf.reg15_q\[26\] _03373_ _03374_ u_rf.reg24_q\[26\] _03905_ VGND VGND VPWR
+ VPWR _03906_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_1_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ u_rf.reg9_q\[23\] _03293_ _03349_ u_rf.reg20_q\[23\] VGND VGND VPWR VPWR
+ _03840_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11670_ _05700_ _02306_ _05709_ VGND VGND VPWR VPWR _01037_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10621_ _05153_ VGND VGND VPWR VPWR _00544_ sky130_fd_sc_hd__clkbuf_1
X_10552_ u_rf.reg16_q\[0\] _04935_ _05116_ VGND VGND VPWR VPWR _05117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10483_ _05079_ VGND VGND VPWR VPWR _00480_ sky130_fd_sc_hd__clkbuf_1
X_12222_ clknet_leaf_12_clk _00259_ net243 VGND VGND VPWR VPWR u_rf.reg8_q\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12153_ clknet_leaf_58_clk _00190_ net291 VGND VGND VPWR VPWR u_rf.reg5_q\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12084_ clknet_leaf_33_clk _00121_ net269 VGND VGND VPWR VPWR u_rf.reg3_q\[25\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11104_ _05409_ VGND VGND VPWR VPWR _00771_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11035_ _04728_ u_rf.reg23_q\[3\] _05369_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ clknet_leaf_94_clk _01023_ net340 VGND VGND VPWR VPWR u_rf.reg31_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11937_ clknet_leaf_74_clk u_decod.rs1_data\[25\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11868_ clknet_leaf_60_clk _00095_ net340 VGND VGND VPWR VPWR u_rf.reg0_q\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11799_ clknet_leaf_76_clk net152 net369 VGND VGND VPWR VPWR u_decod.pc0_q_i\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10819_ _05257_ VGND VGND VPWR VPWR _00638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06010_ u_decod.rs2_data_q\[27\] u_decod.rs1_data_q\[27\] VGND VGND VPWR VPWR _01281_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07961_ _03167_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[32\] sky130_fd_sc_hd__clkbuf_1
X_09700_ _04629_ VGND VGND VPWR VPWR _00147_ sky130_fd_sc_hd__clkbuf_1
X_06912_ u_rf.reg0_q\[10\] _01516_ _01599_ u_rf.reg15_q\[10\] _02161_ VGND VGND VPWR
+ VPWR _02162_ sky130_fd_sc_hd__a221o_1
X_07892_ _02334_ _03086_ _03087_ _03102_ VGND VGND VPWR VPWR _03103_ sky130_fd_sc_hd__o31a_1
XFILLER_0_156_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09631_ _04592_ VGND VGND VPWR VPWR _00115_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06843_ u_decod.rs2_data_q\[0\] _02095_ _01504_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__o21a_1
X_09562_ _04532_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__clkbuf_8
X_06774_ u_rf.reg13_q\[7\] _01597_ _01605_ u_rf.reg3_q\[7\] _02029_ VGND VGND VPWR
+ VPWR _02030_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08513_ u_rf.reg1_q\[16\] _03311_ _03313_ u_rf.reg14_q\[16\] _03700_ VGND VGND VPWR
+ VPWR _03701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09493_ _04495_ VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__buf_6
XFILLER_0_78_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08444_ _03628_ _03630_ _03632_ _03634_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08375_ u_rf.reg8_q\[10\] _03271_ _03273_ u_rf.reg29_q\[10\] _03568_ VGND VGND VPWR
+ VPWR _03569_ sky130_fd_sc_hd__a221o_1
X_07326_ _02553_ _02555_ _02557_ _02559_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07257_ _02288_ _02493_ _01472_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07188_ _02423_ _02425_ _02427_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__or3_1
X_06208_ _01478_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__buf_2
X_06139_ u_decod.rs2_data_q\[25\] u_decod.rs1_data_q\[25\] VGND VGND VPWR VPWR _01410_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_72_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ u_rf.reg6_q\[14\] _04457_ _04695_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__mux2_1
X_12840_ clknet_leaf_21_clk _00877_ net286 VGND VGND VPWR VPWR u_rf.reg27_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_87_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_223 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_109_clk _00808_ net313 VGND VGND VPWR VPWR u_rf.reg25_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11722_ clknet_leaf_25_clk _00014_ net265 VGND VGND VPWR VPWR u_rf.reg2_q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_289 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11653_ _05693_ u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10604_ u_rf.reg16_q\[25\] _04991_ _05138_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_862 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11584_ _05663_ VGND VGND VPWR VPWR _00997_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10535_ _05106_ VGND VGND VPWR VPWR _00505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10466_ _04774_ u_rf.reg14_q\[25\] _05064_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12205_ clknet_leaf_8_clk _00242_ net217 VGND VGND VPWR VPWR u_rf.reg7_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_10397_ _05033_ VGND VGND VPWR VPWR _00440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12136_ clknet_leaf_18_clk _00173_ net288 VGND VGND VPWR VPWR u_rf.reg5_q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12067_ clknet_leaf_108_clk _00104_ net312 VGND VGND VPWR VPWR u_rf.reg3_q\[8\] sky130_fd_sc_hd__dfrtp_1
X_11018_ _05363_ VGND VGND VPWR VPWR _00731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12969_ clknet_leaf_21_clk _01006_ net282 VGND VGND VPWR VPWR u_rf.reg31_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_138_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_138_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06490_ _01688_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_138_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08160_ u_rf.reg28_q\[1\] _03330_ _03332_ u_rf.reg2_q\[1\] VGND VGND VPWR VPWR _03363_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07111_ net133 _02342_ _02344_ _02353_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08091_ _03213_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__buf_8
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07042_ u_decod.rs1_data_q\[28\] _01446_ _01753_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_41_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ u_decod.rs1_data_q\[26\] u_decod.branch_imm_q_o\[26\] VGND VGND VPWR VPWR
+ _04142_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07944_ _03145_ _03147_ _03149_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__or4_1
XFILLER_0_48_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07875_ u_decod.pc_q_o\[29\] _02999_ u_decod.pc_q_o\[30\] VGND VGND VPWR VPWR _03086_
+ sky130_fd_sc_hd__a21oi_1
X_06826_ u_rf.reg23_q\[8\] _01611_ _01655_ u_rf.reg10_q\[8\] _02079_ VGND VGND VPWR
+ VPWR _02080_ sky130_fd_sc_hd__a221o_1
X_09614_ u_rf.reg3_q\[11\] _04451_ _04582_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_129_clk sky130_fd_sc_hd__clkbuf_16
X_09545_ _04546_ VGND VGND VPWR VPWR _00075_ sky130_fd_sc_hd__clkbuf_1
X_06757_ _02013_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[7\] sky130_fd_sc_hd__inv_2
XFILLER_0_78_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06688_ _01311_ _01860_ _01333_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__o21a_1
X_09476_ _04509_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08427_ u_rf.reg7_q\[12\] _03428_ _03429_ u_rf.reg25_q\[12\] _03618_ VGND VGND VPWR
+ VPWR _03619_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08358_ u_rf.reg7_q\[9\] _03369_ _03370_ u_rf.reg25_q\[9\] _03552_ VGND VGND VPWR
+ VPWR _03553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08289_ _03482_ _03484_ _03486_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__or3_1
X_07309_ _02189_ _02543_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10320_ u_decod.rf_ff_res_data_i\[24\] VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10251_ _04942_ VGND VGND VPWR VPWR _00385_ sky130_fd_sc_hd__clkbuf_1
X_10182_ _04728_ u_rf.reg11_q\[3\] _04900_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__mux2_1
Xfanout250 net252 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_4
Xfanout272 net273 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__buf_2
Xfanout261 net264 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout283 net310 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__buf_2
Xfanout294 net297 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_4
X_12823_ clknet_leaf_72_clk _00860_ net359 VGND VGND VPWR VPWR u_rf.reg26_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12754_ clknet_leaf_39_clk _00791_ net277 VGND VGND VPWR VPWR u_rf.reg24_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11705_ _05727_ VGND VGND VPWR VPWR _01054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12685_ clknet_leaf_7_clk _00722_ net218 VGND VGND VPWR VPWR u_rf.reg22_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11636_ _05690_ VGND VGND VPWR VPWR _01022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_507 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11567_ _04784_ u_rf.reg30_q\[30\] _05620_ VGND VGND VPWR VPWR _05654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10518_ _05097_ VGND VGND VPWR VPWR _00497_ sky130_fd_sc_hd__clkbuf_1
X_11498_ _05617_ VGND VGND VPWR VPWR _00957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10449_ _04757_ u_rf.reg14_q\[17\] _05053_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12119_ clknet_leaf_71_clk _00156_ net358 VGND VGND VPWR VPWR u_rf.reg4_q\[28\] sky130_fd_sc_hd__dfrtp_1
X_05990_ u_decod.rs2_data_q\[29\] u_decod.rs1_data_q\[29\] VGND VGND VPWR VPWR _01261_
+ sky130_fd_sc_hd__nor2_1
X_07660_ _02618_ _02880_ _01057_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__a21o_1
X_07591_ _02813_ _02814_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[23\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06611_ _01873_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[4\] sky130_fd_sc_hd__inv_2
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _04409_ u_decod.rs2_data_q\[26\] _04410_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06542_ _01463_ _01806_ _01451_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__mux2_1
X_09261_ _04362_ _04365_ _04366_ _04369_ _04368_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__a41o_1
XFILLER_0_8_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06473_ _01197_ _01232_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__nor2_1
X_08212_ u_rf.reg4_q\[3\] _03356_ _03357_ u_rf.reg17_q\[3\] VGND VGND VPWR VPWR _03413_
+ sky130_fd_sc_hd__a22o_1
X_09192_ _04307_ _04314_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08143_ u_rf.reg26_q\[1\] _03344_ _03345_ u_rf.reg21_q\[1\] VGND VGND VPWR VPWR _03346_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08074_ u_rf.reg22_q\[0\] _03275_ _03277_ u_rf.reg3_q\[0\] VGND VGND VPWR VPWR _03278_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07025_ u_rf.reg1_q\[12\] _01586_ _01666_ u_rf.reg8_q\[12\] VGND VGND VPWR VPWR _02271_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08976_ _04126_ _04127_ VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__xnor2_1
Xhold69 u_decod.pc0_q_i\[21\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _02874_ _02964_ _03051_ _03135_ _01477_ _02685_ VGND VGND VPWR VPWR _03136_
+ sky130_fd_sc_hd__mux4_1
X_07858_ u_rf.reg28_q\[29\] _02419_ _02360_ u_rf.reg9_q\[29\] VGND VGND VPWR VPWR
+ _03070_ sky130_fd_sc_hd__a22o_1
X_07789_ _01266_ _03003_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06809_ _02063_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[8\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09528_ _04537_ VGND VGND VPWR VPWR _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _04500_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__clkbuf_1
X_12470_ clknet_leaf_49_clk _00507_ net306 VGND VGND VPWR VPWR u_rf.reg15_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11421_ u_rf.reg28_q\[25\] u_decod.rf_ff_res_data_i\[25\] _05571_ VGND VGND VPWR
+ VPWR _05577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11352_ _05540_ VGND VGND VPWR VPWR _00888_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_115_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10303_ _04977_ VGND VGND VPWR VPWR _00402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11283_ u_rf.reg26_q\[24\] net477 _05499_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__mux2_1
X_10234_ _04780_ u_rf.reg11_q\[28\] _04922_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__mux2_1
X_10165_ u_rf.reg10_q\[28\] _04486_ _04885_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__mux2_1
X_10096_ _04857_ VGND VGND VPWR VPWR _00315_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12806_ clknet_leaf_3_clk _00843_ net213 VGND VGND VPWR VPWR u_rf.reg26_q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10998_ u_rf.reg22_q\[18\] _04976_ _05344_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_106_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12737_ clknet_leaf_117_clk _00774_ net325 VGND VGND VPWR VPWR u_rf.reg24_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ clknet_leaf_127_clk _00705_ net235 VGND VGND VPWR VPWR u_rf.reg22_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11619_ _04768_ u_rf.reg31_q\[22\] _05679_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12599_ clknet_leaf_70_clk _00636_ net353 VGND VGND VPWR VPWR u_rf.reg19_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_115_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08830_ _04001_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_146_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ u_rf.reg8_q\[28\] _03407_ _03408_ u_rf.reg29_q\[28\] _03936_ VGND VGND VPWR
+ VPWR _03937_ sky130_fd_sc_hd__a221o_1
X_05973_ _01239_ _01090_ _01198_ VGND VGND VPWR VPWR _01249_ sky130_fd_sc_hd__o21a_1
X_08692_ u_rf.reg7_q\[24\] _03428_ _03429_ u_rf.reg25_q\[24\] _03871_ VGND VGND VPWR
+ VPWR _03872_ sky130_fd_sc_hd__a221o_1
X_07712_ u_decod.dec0.funct7\[1\] _01224_ _02646_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__a21o_2
X_07643_ net199 _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07574_ u_rf.reg11_q\[23\] _02375_ _01668_ u_rf.reg8_q\[23\] _02797_ VGND VGND VPWR
+ VPWR _02798_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_124_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09313_ _04404_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_2
X_06525_ _01656_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09244_ _04357_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_62_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06456_ u_rf.reg13_q\[1\] _01597_ _01641_ u_rf.reg26_q\[1\] VGND VGND VPWR VPWR _01724_
+ sky130_fd_sc_hd__a22o_1
X_09175_ u_decod.pc_q_o\[17\] u_decod.branch_imm_q_o\[17\] VGND VGND VPWR VPWR _04300_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_618 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08126_ _03242_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06387_ _01512_ _01553_ _01577_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__and3_2
XFILLER_0_114_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_133_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08057_ _03197_ VGND VGND VPWR VPWR _03261_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07008_ _02233_ _02242_ _02254_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_110_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08959_ _01358_ u_decod.branch_imm_q_o\[21\] VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__xor2_1
X_11970_ clknet_leaf_79_clk net454 net372 VGND VGND VPWR VPWR u_decod.pc_q_o\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_10921_ _05312_ VGND VGND VPWR VPWR _00685_ sky130_fd_sc_hd__clkbuf_1
X_10852_ _05275_ VGND VGND VPWR VPWR _00653_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10783_ u_rf.reg19_q\[13\] _04966_ _05235_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_51_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12522_ clknet_leaf_30_clk _00559_ net261 VGND VGND VPWR VPWR u_rf.reg17_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_229 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ clknet_leaf_121_clk _00490_ net247 VGND VGND VPWR VPWR u_rf.reg15_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_10_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11404_ u_rf.reg28_q\[17\] u_decod.rf_ff_res_data_i\[17\] _05560_ VGND VGND VPWR
+ VPWR _05568_ sky130_fd_sc_hd__mux2_1
X_12384_ clknet_leaf_115_clk _00421_ net323 VGND VGND VPWR VPWR u_rf.reg13_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11335_ _05531_ VGND VGND VPWR VPWR _00880_ sky130_fd_sc_hd__clkbuf_1
X_11266_ u_rf.reg26_q\[16\] u_decod.rf_ff_res_data_i\[16\] _05488_ VGND VGND VPWR
+ VPWR _05495_ sky130_fd_sc_hd__mux2_1
X_13005_ clknet_leaf_65_clk _01042_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[18\]
+ sky130_fd_sc_hd__dfxtp_2
X_10217_ _04899_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11197_ _05458_ VGND VGND VPWR VPWR _00815_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10148_ _04862_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10079_ _04848_ VGND VGND VPWR VPWR _00307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07290_ u_rf.reg17_q\[17\] _01630_ _01656_ u_rf.reg10_q\[17\] _02525_ VGND VGND VPWR
+ VPWR _02526_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06310_ _01579_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__buf_8
XFILLER_0_45_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06241_ _01511_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06172_ _01442_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09931_ _04721_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09862_ u_rf.reg6_q\[30\] _04490_ _04683_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__mux2_1
X_08813_ u_rf.reg0_q\[30\] _03175_ _03241_ u_rf.reg12_q\[30\] _03986_ VGND VGND VPWR
+ VPWR _03987_ sky130_fd_sc_hd__a221o_1
X_09793_ u_rf.reg5_q\[30\] _04490_ _04646_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__mux2_1
X_08744_ u_rf.reg31_q\[27\] _03504_ _03505_ u_rf.reg11_q\[27\] _03920_ VGND VGND VPWR
+ VPWR _03921_ sky130_fd_sc_hd__a221o_1
X_05956_ _01231_ _01085_ _01209_ _01235_ VGND VGND VPWR VPWR _01236_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05887_ net484 _01142_ _01119_ net83 _01182_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__a221o_1
X_08675_ net439 _03773_ _03855_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07626_ u_rf.reg25_q\[24\] _01783_ _02367_ u_rf.reg14_q\[24\] VGND VGND VPWR VPWR
+ _02848_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07557_ _01368_ _01820_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_33_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
X_06508_ u_decod.dec0.instr_i\[9\] _01226_ _01715_ u_decod.dec0.instr_i\[22\] VGND
+ VGND VPWR VPWR _01774_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07488_ _02699_ _02706_ _02715_ _01680_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__o31a_2
XFILLER_0_91_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09227_ _04136_ _04206_ _04275_ _04344_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[24\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06439_ _01503_ _01707_ _01478_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_267 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09158_ _04279_ _04272_ _04276_ _04277_ _04285_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_79_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08109_ _03312_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__buf_8
X_09089_ u_decod.pc_q_o\[5\] u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _04226_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11120_ u_rf.reg24_q\[11\] _04962_ _05416_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11051_ _05381_ VGND VGND VPWR VPWR _00746_ sky130_fd_sc_hd__clkbuf_1
X_10002_ _04807_ VGND VGND VPWR VPWR _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11953_ clknet_leaf_100_clk net391 net338 VGND VGND VPWR VPWR u_decod.pc_q_o\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_123_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10904_ _05303_ VGND VGND VPWR VPWR _00677_ sky130_fd_sc_hd__clkbuf_1
X_11884_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[5\] net322 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10835_ _05266_ VGND VGND VPWR VPWR _00645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10766_ u_rf.reg19_q\[5\] _04949_ _05224_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12505_ clknet_leaf_58_clk _00542_ net292 VGND VGND VPWR VPWR u_rf.reg16_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10697_ _05193_ VGND VGND VPWR VPWR _00580_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12436_ clknet_leaf_31_clk _00473_ net261 VGND VGND VPWR VPWR u_rf.reg14_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_187 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12367_ clknet_leaf_42_clk _00404_ net276 VGND VGND VPWR VPWR u_rf.reg12_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12298_ clknet_leaf_30_clk _00335_ net261 VGND VGND VPWR VPWR u_rf.reg10_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11318_ _05522_ VGND VGND VPWR VPWR _00872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11249_ u_rf.reg26_q\[8\] u_decod.rf_ff_res_data_i\[8\] _05477_ VGND VGND VPWR VPWR
+ _05486_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05810_ u_decod.pc0_q_i\[6\] u_decod.pc0_q_i\[7\] u_decod.pc0_q_i\[8\] _01113_ VGND
+ VGND VPWR VPWR _01124_ sky130_fd_sc_hd__and4_1
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06790_ _01957_ _02044_ _01474_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__mux2_1
X_05741_ _01062_ _01065_ VGND VGND VPWR VPWR _01066_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08460_ u_rf.reg31_q\[14\] _03210_ _03291_ u_rf.reg11_q\[14\] VGND VGND VPWR VPWR
+ _03650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07411_ _02622_ _02634_ _02641_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__or3b_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08391_ u_decod.exe_ff_res_data_i\[10\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[10\]
+ _03584_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07342_ _01386_ _02534_ _01379_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_15_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07273_ u_decod.dec0.instr_i\[17\] _01208_ _02256_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__a21o_1
XFILLER_0_73_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_154_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09012_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__and2b_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06224_ _01061_ _01445_ _01494_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_154_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold100 u_decod.pc0_q_i\[8\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06155_ _01061_ _01425_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold133 u_exe.pc_data_q\[13\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 u_decod.branch_imm_q_o\[14\] VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 u_decod.dec0.funct7\[4\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 u_decod.rf_ff_res_data_i\[1\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_1
Xhold155 u_rf.reg16_q\[29\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06086_ _01290_ _01294_ _01356_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_57_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09914_ _04752_ VGND VGND VPWR VPWR _00238_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09845_ _04708_ VGND VGND VPWR VPWR _00213_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09776_ _04671_ VGND VGND VPWR VPWR _00181_ sky130_fd_sc_hd__clkbuf_1
X_06988_ u_decod.pc_q_o\[12\] _02185_ _01484_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__o21ai_1
X_08727_ u_rf.reg6_q\[26\] _03304_ _03306_ u_rf.reg13_q\[26\] VGND VGND VPWR VPWR
+ _03905_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05939_ _01071_ _01086_ _01084_ _01221_ VGND VGND VPWR VPWR _01222_ sky130_fd_sc_hd__and4_1
X_08658_ u_rf.reg18_q\[23\] _03353_ _03355_ u_rf.reg23_q\[23\] _03838_ VGND VGND VPWR
+ VPWR _03839_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_438 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ net49 net100 _02446_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__a21bo_1
X_08589_ _03257_ VGND VGND VPWR VPWR _03773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10620_ u_rf.reg17_q\[0\] _04935_ _05152_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_335 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10551_ _05115_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10482_ _04719_ u_rf.reg15_q\[0\] _05078_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_278 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12221_ clknet_leaf_16_clk _00258_ net250 VGND VGND VPWR VPWR u_rf.reg8_q\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12152_ clknet_leaf_66_clk _00189_ net349 VGND VGND VPWR VPWR u_rf.reg5_q\[29\] sky130_fd_sc_hd__dfrtp_1
X_12083_ clknet_leaf_51_clk _00120_ net304 VGND VGND VPWR VPWR u_rf.reg3_q\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11103_ u_rf.reg24_q\[3\] _04945_ _05405_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__mux2_1
X_11034_ _05372_ VGND VGND VPWR VPWR _00738_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ clknet_leaf_64_clk _01022_ net346 VGND VGND VPWR VPWR u_rf.reg31_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_11936_ clknet_leaf_74_clk u_decod.rs1_data\[24\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11867_ clknet_leaf_57_clk _00094_ net343 VGND VGND VPWR VPWR u_rf.reg0_q\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ clknet_leaf_80_clk net151 net370 VGND VGND VPWR VPWR u_decod.pc0_q_i\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10818_ u_rf.reg19_q\[30\] _05001_ _05223_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10749_ _05220_ VGND VGND VPWR VPWR _00605_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12419_ clknet_leaf_108_clk _00456_ net312 VGND VGND VPWR VPWR u_rf.reg14_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07960_ _03165_ _03166_ _03164_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_06911_ u_rf.reg7_q\[10\] _01559_ _01604_ u_rf.reg3_q\[10\] VGND VGND VPWR VPWR _02161_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07891_ _03088_ _03094_ _03096_ _03098_ _03101_ VGND VGND VPWR VPWR _03102_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09630_ u_rf.reg3_q\[19\] _04467_ _04582_ VGND VGND VPWR VPWR _04592_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06842_ _01824_ _01904_ _02001_ _02094_ _01474_ _01458_ VGND VGND VPWR VPWR _02095_
+ sky130_fd_sc_hd__mux4_2
X_09561_ _04554_ VGND VGND VPWR VPWR _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06773_ u_rf.reg7_q\[7\] _01559_ _01672_ u_rf.reg2_q\[7\] VGND VGND VPWR VPWR _02029_
+ sky130_fd_sc_hd__a22o_1
X_08512_ u_rf.reg7_q\[16\] _03314_ _03315_ u_rf.reg25_q\[16\] VGND VGND VPWR VPWR
+ _03700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09492_ _04517_ VGND VGND VPWR VPWR _00051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08443_ u_rf.reg26_q\[13\] _03344_ _03357_ u_rf.reg17_q\[13\] _03633_ VGND VGND VPWR
+ VPWR _03634_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08374_ u_rf.reg22_q\[10\] _03275_ _03277_ u_rf.reg3_q\[10\] VGND VGND VPWR VPWR
+ _03568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07325_ u_rf.reg31_q\[18\] _01616_ _01659_ u_rf.reg14_q\[18\] _02558_ VGND VGND VPWR
+ VPWR _02559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07256_ _01468_ _02099_ _01498_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__o21a_1
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_647 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06207_ u_decod.rs2_data_q\[0\] VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__inv_2
XFILLER_0_131_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07187_ u_rf.reg0_q\[15\] _01664_ _02360_ u_rf.reg9_q\[15\] _02426_ VGND VGND VPWR
+ VPWR _02427_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06138_ u_decod.rs2_data_q\[26\] u_decod.rs1_data_q\[26\] VGND VGND VPWR VPWR _01409_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06069_ _01338_ _01339_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_107_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _04699_ VGND VGND VPWR VPWR _00205_ sky130_fd_sc_hd__clkbuf_1
X_09759_ _04662_ VGND VGND VPWR VPWR _00173_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12770_ clknet_leaf_127_clk _00807_ net235 VGND VGND VPWR VPWR u_rf.reg25_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11721_ clknet_leaf_19_clk _00013_ net281 VGND VGND VPWR VPWR u_rf.reg2_q\[13\] sky130_fd_sc_hd__dfrtp_1
X_11652_ net345 VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _05143_ VGND VGND VPWR VPWR _00536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11583_ _04732_ u_rf.reg31_q\[5\] _05657_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10534_ _04774_ u_rf.reg15_q\[25\] _05100_ VGND VGND VPWR VPWR _05106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10465_ _05069_ VGND VGND VPWR VPWR _00472_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10396_ _04772_ u_rf.reg13_q\[24\] _05028_ VGND VGND VPWR VPWR _05033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12204_ clknet_leaf_19_clk _00241_ net281 VGND VGND VPWR VPWR u_rf.reg7_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12135_ clknet_leaf_4_clk _00172_ net211 VGND VGND VPWR VPWR u_rf.reg5_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_12066_ clknet_leaf_131_clk _00103_ net229 VGND VGND VPWR VPWR u_rf.reg3_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11017_ u_rf.reg22_q\[27\] _04995_ _05355_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12968_ clknet_leaf_17_clk _01005_ net289 VGND VGND VPWR VPWR u_rf.reg31_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12899_ clknet_leaf_108_clk _00936_ net314 VGND VGND VPWR VPWR u_rf.reg29_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11919_ clknet_leaf_102_clk u_decod.rs1_data\[7\] net337 VGND VGND VPWR VPWR u_decod.rs1_data_q\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_138_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07110_ _01425_ _02290_ _02352_ _01442_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08090_ _03293_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07041_ u_decod.rs1_data_q\[20\] _01454_ _01753_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ _04101_ _04141_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_54_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07943_ u_rf.reg31_q\[31\] _01777_ _02380_ u_rf.reg10_q\[31\] _03150_ VGND VGND VPWR
+ VPWR _03151_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07874_ _01273_ _03083_ _01765_ VGND VGND VPWR VPWR _03085_ sky130_fd_sc_hd__a21o_1
X_06825_ u_rf.reg6_q\[8\] _01554_ _01651_ u_rf.reg22_q\[8\] VGND VGND VPWR VPWR _02079_
+ sky130_fd_sc_hd__a22o_1
X_09613_ _04583_ VGND VGND VPWR VPWR _00106_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09544_ u_rf.reg0_q\[11\] _04451_ _04544_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__mux2_1
X_06756_ _01765_ _01993_ _01998_ _02004_ _02012_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09475_ u_rf.reg1_q\[11\] _04451_ _04507_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__mux2_1
X_06687_ _01944_ _01946_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[5\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08426_ u_rf.reg1_q\[12\] _03446_ _03447_ u_rf.reg14_q\[12\] VGND VGND VPWR VPWR
+ _03618_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_498 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_329 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_148 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08357_ u_rf.reg1_q\[9\] _03310_ _03312_ u_rf.reg14_q\[9\] VGND VGND VPWR VPWR _03552_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08288_ u_rf.reg27_q\[6\] _03318_ _03320_ u_rf.reg19_q\[6\] _03485_ VGND VGND VPWR
+ VPWR _03486_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07308_ _01475_ _02450_ _02542_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07239_ u_rf.reg23_q\[16\] _01612_ _01621_ u_rf.reg24_q\[16\] VGND VGND VPWR VPWR
+ _02477_ sky130_fd_sc_hd__a22o_1
X_10250_ u_rf.reg12_q\[1\] _04941_ _04939_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10181_ _04903_ VGND VGND VPWR VPWR _00354_ sky130_fd_sc_hd__clkbuf_1
Xfanout240 net254 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__buf_2
Xfanout273 net274 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_4
Xfanout262 net264 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout251 net252 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_4
Xfanout295 net297 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_2
Xfanout284 net287 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_4
X_12822_ clknet_leaf_72_clk _00859_ net358 VGND VGND VPWR VPWR u_rf.reg26_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12753_ clknet_leaf_21_clk _00790_ net286 VGND VGND VPWR VPWR u_rf.reg24_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11704_ u_decod.branch_imm_q_o\[30\] _03105_ _05717_ VGND VGND VPWR VPWR _05727_
+ sky130_fd_sc_hd__mux2_1
X_12684_ clknet_leaf_26_clk _00721_ net265 VGND VGND VPWR VPWR u_rf.reg22_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11635_ _04784_ u_rf.reg31_q\[30\] _05656_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11566_ _05653_ VGND VGND VPWR VPWR _00989_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_519 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10517_ _04757_ u_rf.reg15_q\[17\] _05089_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11497_ _04782_ u_rf.reg29_q\[29\] _05607_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__mux2_1
X_10448_ _05060_ VGND VGND VPWR VPWR _00464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10379_ _04755_ u_rf.reg13_q\[16\] _05017_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12118_ clknet_leaf_51_clk _00155_ net308 VGND VGND VPWR VPWR u_rf.reg4_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_396 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12049_ clknet_leaf_65_clk u_decod.exe_ff_res_data_i\[29\] net357 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[29\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07590_ net200 _02768_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__nor2_1
X_06610_ net133 _01856_ _01863_ _01872_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__a211oi_2
X_06541_ _01384_ _01683_ _01302_ u_decod.rs1_data_q\[26\] _01446_ _01685_ VGND VGND
+ VPWR VPWR _01806_ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09260_ u_decod.pc_q_o\[29\] u_decod.branch_imm_q_o\[29\] VGND VGND VPWR VPWR _04373_
+ sky130_fd_sc_hd__and2_1
X_06472_ u_decod.dec0.funct7\[3\] u_decod.dec0.funct7\[2\] u_decod.dec0.funct7\[4\]
+ _01081_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__nor4_1
XFILLER_0_146_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08211_ u_rf.reg8_q\[3\] _03407_ _03408_ u_rf.reg29_q\[3\] _03411_ VGND VGND VPWR
+ VPWR _03412_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09191_ _04296_ _04303_ _04301_ _04308_ _04300_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a311o_1
XFILLER_0_90_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08142_ _03285_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08073_ _03276_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__buf_8
XFILLER_0_43_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07024_ u_rf.reg17_q\[12\] _01631_ _01791_ u_rf.reg10_q\[12\] _02269_ VGND VGND VPWR
+ VPWR _02270_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08975_ _04119_ _04122_ _04117_ VGND VGND VPWR VPWR _04127_ sky130_fd_sc_hd__o21a_1
X_07926_ _01267_ _01367_ _01289_ u_decod.rs1_data_q\[7\] _01469_ _01466_ VGND VGND
+ VPWR VPWR _03135_ sky130_fd_sc_hd__mux4_1
X_07857_ _03062_ _03064_ _03066_ _03068_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__or4_1
X_07788_ _01287_ _03002_ _01413_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06808_ _01441_ _02041_ _02062_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06739_ _01910_ _01995_ _01315_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__mux2_1
X_09527_ u_rf.reg0_q\[3\] _04434_ _04533_ VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09458_ u_rf.reg1_q\[3\] _04434_ _04496_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09389_ u_rf.reg2_q\[12\] _04453_ _04449_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__mux2_1
X_08409_ u_rf.reg28_q\[11\] _03331_ _03333_ u_rf.reg2_q\[11\] VGND VGND VPWR VPWR
+ _03602_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11420_ _05576_ VGND VGND VPWR VPWR _00920_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11351_ _04772_ u_rf.reg27_q\[24\] _05535_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_115_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10302_ u_rf.reg12_q\[18\] _04976_ _04960_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__mux2_1
X_11282_ _05503_ VGND VGND VPWR VPWR _00855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10233_ _04930_ VGND VGND VPWR VPWR _00379_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10164_ _04893_ VGND VGND VPWR VPWR _00347_ sky130_fd_sc_hd__clkbuf_1
X_10095_ u_rf.reg9_q\[27\] _04484_ _04849_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12805_ clknet_leaf_116_clk _00842_ net324 VGND VGND VPWR VPWR u_rf.reg26_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10997_ _05352_ VGND VGND VPWR VPWR _00721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12736_ clknet_leaf_116_clk _00773_ net327 VGND VGND VPWR VPWR u_rf.reg24_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12667_ clknet_leaf_11_clk _00704_ net222 VGND VGND VPWR VPWR u_rf.reg22_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11618_ _05681_ VGND VGND VPWR VPWR _01013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12598_ clknet_leaf_47_clk _00635_ net306 VGND VGND VPWR VPWR u_rf.reg19_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11549_ _04766_ u_rf.reg30_q\[21\] _05643_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_146_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ u_rf.reg22_q\[28\] _03274_ _03276_ u_rf.reg3_q\[28\] VGND VGND VPWR VPWR
+ _03936_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05972_ _01224_ _01222_ VGND VGND VPWR VPWR _01248_ sky130_fd_sc_hd__or2_1
X_07711_ _02929_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[26\] sky130_fd_sc_hd__inv_2
X_08691_ u_rf.reg1_q\[24\] _03311_ _03313_ u_rf.reg14_q\[24\] VGND VGND VPWR VPWR
+ _03871_ sky130_fd_sc_hd__a22o_1
X_07642_ _02089_ _02487_ _02863_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_49_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07573_ u_rf.reg6_q\[23\] _01557_ _01653_ u_rf.reg22_q\[23\] VGND VGND VPWR VPWR
+ _02797_ sky130_fd_sc_hd__a22o_1
X_09312_ _04397_ u_decod.rs2_data_q\[18\] _04398_ VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06524_ _01782_ _01786_ _01789_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__or3_1
XFILLER_0_146_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09243_ _04351_ _04353_ _04350_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_76_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06455_ u_rf.reg5_q\[1\] _01568_ _01666_ u_rf.reg8_q\[1\] _01722_ VGND VGND VPWR
+ VPWR _01723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09174_ _04090_ _04274_ _04275_ _04299_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[16\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_282 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06386_ _01655_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_32_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08125_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08056_ _03187_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__buf_2
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07007_ _01059_ _02243_ _02246_ _02253_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08958_ _04101_ _04112_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__nor2_1
X_07909_ u_rf.reg23_q\[30\] _02652_ _02385_ u_rf.reg20_q\[30\] VGND VGND VPWR VPWR
+ _03119_ sky130_fd_sc_hd__a22o_1
X_08889_ _04050_ net388 VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__xnor2_1
X_10920_ u_rf.reg21_q\[13\] _04966_ _05308_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10851_ u_rf.reg20_q\[13\] _04966_ _05271_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10782_ _05238_ VGND VGND VPWR VPWR _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12521_ clknet_leaf_23_clk _00558_ net267 VGND VGND VPWR VPWR u_rf.reg17_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ clknet_leaf_111_clk _00489_ net316 VGND VGND VPWR VPWR u_rf.reg15_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11403_ _05567_ VGND VGND VPWR VPWR _00912_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12383_ clknet_leaf_137_clk _00420_ net205 VGND VGND VPWR VPWR u_rf.reg13_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11334_ _04755_ u_rf.reg27_q\[16\] _05524_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__mux2_1
X_11265_ _05494_ VGND VGND VPWR VPWR _00847_ sky130_fd_sc_hd__clkbuf_1
X_13004_ clknet_leaf_65_clk _01041_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[17\]
+ sky130_fd_sc_hd__dfxtp_2
X_10216_ _04921_ VGND VGND VPWR VPWR _00371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11196_ u_rf.reg25_q\[15\] _04970_ _05452_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10147_ _04884_ VGND VGND VPWR VPWR _00339_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10078_ u_rf.reg9_q\[19\] _04467_ _04838_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ clknet_leaf_42_clk _00756_ net275 VGND VGND VPWR VPWR u_rf.reg23_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06240_ _01260_ _01440_ _01510_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_44_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_414 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06171_ _01441_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__buf_2
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09930_ u_decod.rf_ff_res_data_i\[20\] VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09861_ _04716_ VGND VGND VPWR VPWR _00221_ sky130_fd_sc_hd__clkbuf_1
X_09792_ _04679_ VGND VGND VPWR VPWR _00189_ sky130_fd_sc_hd__clkbuf_1
X_08812_ u_rf.reg28_q\[30\] _03242_ _03243_ u_rf.reg2_q\[30\] VGND VGND VPWR VPWR
+ _03986_ sky130_fd_sc_hd__a22o_1
X_08743_ u_rf.reg9_q\[27\] _03293_ _03295_ u_rf.reg20_q\[27\] VGND VGND VPWR VPWR
+ _03920_ sky130_fd_sc_hd__a22o_1
X_05955_ _01080_ _01234_ u_decod.dec0.funct7\[6\] VGND VGND VPWR VPWR _01235_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08674_ u_decod.exe_ff_res_data_i\[23\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[23\]
+ _03854_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__a221o_1
X_05886_ _01180_ _01144_ _01181_ VGND VGND VPWR VPWR _01182_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_37_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ u_rf.reg11_q\[24\] _02375_ _02665_ u_rf.reg19_q\[24\] _02846_ VGND VGND VPWR
+ VPWR _02847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ u_decod.instr_operation_q\[1\] VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__buf_4
XFILLER_0_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06507_ _01714_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__clkbuf_4
X_09226_ _04342_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__xor2_1
X_07487_ _02708_ _02710_ _02712_ _02714_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__or4_1
XFILLER_0_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06438_ _01493_ _01706_ _01502_ VGND VGND VPWR VPWR _01707_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06369_ _01638_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__buf_6
X_09157_ _04276_ u_decod.branch_imm_q_o\[12\] u_decod.pc_q_o\[12\] VGND VGND VPWR
+ VPWR _04285_ sky130_fd_sc_hd__nand3b_1
XTAP_TAPCELL_ROW_79_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08108_ _03232_ VGND VGND VPWR VPWR _03312_ sky130_fd_sc_hd__buf_8
X_09088_ _04017_ _04207_ _04208_ _04225_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[4\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_141_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08039_ u_rf.reg0_q\[31\] _03174_ _03241_ u_rf.reg12_q\[31\] _03244_ VGND VGND VPWR
+ VPWR _03245_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11050_ _04742_ u_rf.reg23_q\[10\] _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__mux2_1
X_10001_ u_rf.reg8_q\[15\] _04459_ _04801_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11952_ clknet_leaf_102_clk net441 net336 VGND VGND VPWR VPWR u_decod.pc_q_o\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10903_ u_rf.reg21_q\[5\] _04949_ _05297_ VGND VGND VPWR VPWR _05303_ sky130_fd_sc_hd__mux2_1
X_11883_ clknet_leaf_102_clk u_decod.rs2_data_nxt\[4\] net335 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10834_ u_rf.reg20_q\[5\] _04949_ _05260_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12504_ clknet_leaf_52_clk _00541_ net304 VGND VGND VPWR VPWR u_rf.reg16_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10765_ _05229_ VGND VGND VPWR VPWR _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10696_ u_rf.reg18_q\[4\] _04947_ _05188_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__mux2_1
X_12435_ clknet_leaf_67_clk _00472_ net350 VGND VGND VPWR VPWR u_rf.reg14_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12366_ clknet_leaf_7_clk _00403_ net216 VGND VGND VPWR VPWR u_rf.reg12_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11317_ _04738_ u_rf.reg27_q\[8\] _05513_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12297_ clknet_leaf_24_clk _00334_ net267 VGND VGND VPWR VPWR u_rf.reg10_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11248_ _05485_ VGND VGND VPWR VPWR _00839_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11179_ u_rf.reg25_q\[7\] _04953_ _05441_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05740_ u_decod.branch_imm_q_o\[0\] _01061_ VGND VGND VPWR VPWR _01065_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07410_ _01765_ _02636_ _02637_ _02640_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o31a_1
X_08390_ _03574_ _03583_ _03337_ VGND VGND VPWR VPWR _03584_ sky130_fd_sc_hd__o21a_1
X_07341_ _02572_ _02574_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[18\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07272_ _01437_ _02490_ _02491_ _02505_ _02508_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[17\]
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09011_ u_decod.rs1_data_q\[28\] u_decod.branch_imm_q_o\[28\] VGND VGND VPWR VPWR
+ _04158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_712 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06223_ u_decod.rs1_data_q\[31\] u_decod.instr_operation_q\[2\] _01445_ VGND VGND
+ VPWR VPWR _01494_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 u_decod.pc0_q_i\[7\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_2
X_06154_ _01424_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__buf_2
XFILLER_0_123_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold123 u_decod.pc0_q_i\[6\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 u_decod.dec0.instr_i\[9\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 u_rf.reg0_q\[25\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__dlygate4sd3_1
X_06085_ _01295_ _01299_ _01351_ _01352_ _01355_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__o311a_1
Xhold145 u_rf.reg18_q\[17\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _04751_ u_rf.reg7_q\[14\] _04743_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ u_rf.reg6_q\[21\] _04472_ _04706_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09775_ u_rf.reg5_q\[21\] _04472_ _04669_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__mux2_1
X_06987_ u_decod.pc_q_o\[12\] _02185_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__and2_1
X_08726_ _03897_ _03899_ _03901_ _03903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__or4_1
X_05938_ u_decod.dec0.funct3\[1\] _01077_ VGND VGND VPWR VPWR _01221_ sky130_fd_sc_hd__nor2_1
X_08657_ u_rf.reg4_q\[23\] _03265_ _03267_ u_rf.reg17_q\[23\] VGND VGND VPWR VPWR
+ _03838_ sky130_fd_sc_hd__a22o_1
X_05869_ u_decod.pc0_q_i\[20\] u_decod.pc0_q_i\[21\] _01159_ u_decod.pc0_q_i\[22\]
+ VGND VGND VPWR VPWR _01169_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _02723_ _02830_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08588_ net454 _03565_ _03772_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[19\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07539_ _02357_ u_decod.exe_ff_res_data_i\[22\] _02764_ VGND VGND VPWR VPWR _02765_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ _04531_ _05114_ VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__nor2_4
XFILLER_0_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09209_ u_decod.pc_q_o\[22\] u_decod.branch_imm_q_o\[22\] VGND VGND VPWR VPWR _04329_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10481_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12220_ clknet_leaf_128_clk _00257_ net236 VGND VGND VPWR VPWR u_rf.reg8_q\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12151_ clknet_leaf_69_clk _00188_ net354 VGND VGND VPWR VPWR u_rf.reg5_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12082_ clknet_leaf_38_clk _00119_ net277 VGND VGND VPWR VPWR u_rf.reg3_q\[23\] sky130_fd_sc_hd__dfrtp_1
X_11102_ _05408_ VGND VGND VPWR VPWR _00770_ sky130_fd_sc_hd__clkbuf_1
X_11033_ _04726_ u_rf.reg23_q\[2\] _05369_ VGND VGND VPWR VPWR _05372_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ clknet_leaf_52_clk _01021_ net351 VGND VGND VPWR VPWR u_rf.reg31_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11935_ clknet_leaf_78_clk u_decod.rs1_data\[23\] net370 VGND VGND VPWR VPWR u_decod.rs1_data_q\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11866_ clknet_leaf_66_clk _00093_ net355 VGND VGND VPWR VPWR u_rf.reg0_q\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11797_ clknet_leaf_77_clk net150 net372 VGND VGND VPWR VPWR u_decod.pc0_q_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10817_ _05256_ VGND VGND VPWR VPWR _00637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10748_ u_rf.reg18_q\[29\] _04999_ _05210_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10679_ _05183_ VGND VGND VPWR VPWR _00572_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12418_ clknet_leaf_130_clk _00455_ net230 VGND VGND VPWR VPWR u_rf.reg14_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12349_ clknet_leaf_15_clk _00386_ net245 VGND VGND VPWR VPWR u_rf.reg12_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06910_ u_rf.reg1_q\[10\] _01585_ _01634_ u_rf.reg9_q\[10\] _02159_ VGND VGND VPWR
+ VPWR _02160_ sky130_fd_sc_hd__a221o_1
X_07890_ _02723_ _03099_ _03100_ _02789_ VGND VGND VPWR VPWR _03101_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_52_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06841_ _01455_ _01704_ _02093_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__a21o_1
X_09560_ u_rf.reg0_q\[19\] _04467_ _04544_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__mux2_1
X_06772_ u_rf.reg6_q\[7\] _01554_ _01630_ u_rf.reg17_q\[7\] _02027_ VGND VGND VPWR
+ VPWR _02028_ sky130_fd_sc_hd__a221o_1
X_09491_ u_rf.reg1_q\[19\] _04467_ _04507_ VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08511_ _03692_ _03694_ _03696_ _03698_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__or4_1
XFILLER_0_148_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08442_ u_rf.reg12_q\[13\] _03241_ _03223_ u_rf.reg23_q\[13\] VGND VGND VPWR VPWR
+ _03633_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08373_ u_rf.reg18_q\[10\] _03262_ _03263_ u_rf.reg23_q\[10\] _03566_ VGND VGND VPWR
+ VPWR _03567_ sky130_fd_sc_hd__a221o_1
X_07324_ u_rf.reg7_q\[18\] _01561_ _01642_ u_rf.reg26_q\[18\] VGND VGND VPWR VPWR
+ _02558_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07255_ net100 net41 _02446_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06206_ _01476_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07186_ u_rf.reg19_q\[15\] _01595_ _01650_ u_rf.reg4_q\[15\] VGND VGND VPWR VPWR
+ _02426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06137_ _01288_ _01407_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06068_ u_decod.rs2_data_q\[8\] u_decod.rs1_data_q\[8\] VGND VGND VPWR VPWR _01339_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ u_rf.reg6_q\[13\] _04455_ _04695_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__mux2_1
X_09758_ u_rf.reg5_q\[13\] _04455_ _04658_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__mux2_1
X_08709_ u_rf.reg15_q\[25\] _03301_ _03303_ u_rf.reg24_q\[25\] _03887_ VGND VGND VPWR
+ VPWR _03888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ u_rf.reg4_q\[14\] _04457_ _04619_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_87_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ clknet_leaf_4_clk _00012_ net211 VGND VGND VPWR VPWR u_rf.reg2_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11651_ _05699_ VGND VGND VPWR VPWR _01028_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_25_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ u_rf.reg16_q\[24\] _04989_ _05138_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11582_ _05662_ VGND VGND VPWR VPWR _00996_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10533_ _05105_ VGND VGND VPWR VPWR _00504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10464_ _04772_ u_rf.reg14_q\[24\] _05064_ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10395_ _05032_ VGND VGND VPWR VPWR _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12203_ clknet_leaf_1_clk _00240_ net221 VGND VGND VPWR VPWR u_rf.reg7_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12134_ clknet_leaf_140_clk _00171_ net202 VGND VGND VPWR VPWR u_rf.reg5_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12065_ clknet_leaf_17_clk _00102_ net251 VGND VGND VPWR VPWR u_rf.reg3_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11016_ _05362_ VGND VGND VPWR VPWR _00730_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12967_ clknet_leaf_2_clk _01004_ net214 VGND VGND VPWR VPWR u_rf.reg31_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11918_ clknet_leaf_97_clk u_decod.rs1_data\[6\] net332 VGND VGND VPWR VPWR u_decod.rs1_data_q\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12898_ clknet_leaf_130_clk _00935_ net229 VGND VGND VPWR VPWR u_rf.reg29_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_138_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11849_ clknet_leaf_4_clk _00076_ net211 VGND VGND VPWR VPWR u_rf.reg0_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07040_ u_decod.pc_q_o\[13\] _02234_ _01484_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08991_ _04139_ _04140_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_54_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07942_ u_rf.reg12_q\[31\] _01610_ _02697_ u_rf.reg4_q\[31\] VGND VGND VPWR VPWR
+ _03150_ sky130_fd_sc_hd__a22o_1
X_07873_ _01273_ _03083_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__nor2_1
X_06824_ u_rf.reg1_q\[8\] _01585_ _01634_ u_rf.reg9_q\[8\] _02077_ VGND VGND VPWR
+ VPWR _02078_ sky130_fd_sc_hd__a221o_1
X_09612_ u_rf.reg3_q\[10\] _04448_ _04582_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__mux2_1
X_09543_ _04545_ VGND VGND VPWR VPWR _00074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06755_ _01764_ _02005_ _02006_ _02009_ _02011_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_102_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09474_ _04508_ VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__clkbuf_1
X_06686_ _01743_ _01945_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__or2_1
X_08425_ u_rf.reg15_q\[12\] _03373_ _03374_ u_rf.reg24_q\[12\] _03616_ VGND VGND VPWR
+ VPWR _03617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _03544_ _03546_ _03548_ _03550_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07307_ _01688_ _02541_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08287_ u_rf.reg16_q\[6\] _03322_ _03324_ u_rf.reg5_q\[6\] VGND VGND VPWR VPWR _03485_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07238_ _02469_ _02471_ _02473_ _02475_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07169_ net39 _02047_ _02049_ net57 _02051_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10180_ _04726_ u_rf.reg11_q\[2\] _04900_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__mux2_1
Xfanout230 net233 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_2
Xfanout241 net253 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_4
Xfanout274 net311 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_4
Xfanout263 net264 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout252 net253 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_2
Xfanout296 net297 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_4
Xfanout285 net287 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_2
X_12821_ clknet_leaf_44_clk _00858_ net297 VGND VGND VPWR VPWR u_rf.reg26_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12752_ clknet_leaf_36_clk _00789_ net271 VGND VGND VPWR VPWR u_rf.reg24_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11703_ _05726_ VGND VGND VPWR VPWR _01053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12683_ clknet_leaf_1_clk _00720_ net209 VGND VGND VPWR VPWR u_rf.reg22_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_11634_ _05689_ VGND VGND VPWR VPWR _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11565_ _04782_ u_rf.reg30_q\[29\] _05643_ VGND VGND VPWR VPWR _05653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11496_ _05616_ VGND VGND VPWR VPWR _00956_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_133_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10516_ _05096_ VGND VGND VPWR VPWR _00496_ sky130_fd_sc_hd__clkbuf_1
X_10447_ _04755_ u_rf.reg14_q\[16\] _05053_ VGND VGND VPWR VPWR _05060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10378_ _05023_ VGND VGND VPWR VPWR _00431_ sky130_fd_sc_hd__clkbuf_1
X_12117_ clknet_leaf_44_clk _00154_ net294 VGND VGND VPWR VPWR u_rf.reg4_q\[26\] sky130_fd_sc_hd__dfrtp_1
X_12048_ clknet_leaf_66_clk u_decod.exe_ff_res_data_i\[28\] net355 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[28\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06540_ _01802_ _01805_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[2\] sky130_fd_sc_hd__xor2_1
XFILLER_0_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06471_ _01085_ _01738_ _01233_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08210_ u_rf.reg22_q\[3\] _03409_ _03410_ u_rf.reg3_q\[3\] VGND VGND VPWR VPWR _03411_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_190 _01747_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09190_ _04311_ _04312_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_64_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08141_ _03343_ VGND VGND VPWR VPWR _03344_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_114_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08072_ _03219_ VGND VGND VPWR VPWR _03276_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07023_ u_rf.reg29_q\[12\] _01627_ _01653_ u_rf.reg22_q\[12\] VGND VGND VPWR VPWR
+ _02269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08974_ _04124_ _04125_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07925_ _02619_ net57 _02618_ VGND VGND VPWR VPWR _03134_ sky130_fd_sc_hd__a21boi_1
X_07856_ u_rf.reg16_q\[29\] _02307_ _02380_ u_rf.reg10_q\[29\] _03067_ VGND VGND VPWR
+ VPWR _03068_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07787_ _01357_ _01393_ _01407_ VGND VGND VPWR VPWR _03002_ sky130_fd_sc_hd__a21oi_1
X_06807_ _01504_ _02046_ _02058_ _02061_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ _04536_ VGND VGND VPWR VPWR _00066_ sky130_fd_sc_hd__clkbuf_1
X_06738_ _01806_ _01994_ _01450_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09457_ _04499_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06669_ u_rf.reg26_q\[5\] _01641_ _01658_ u_rf.reg14_q\[5\] _01928_ VGND VGND VPWR
+ VPWR _01929_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08408_ u_rf.reg27_q\[11\] _03319_ _03321_ u_rf.reg19_q\[11\] _03600_ VGND VGND VPWR
+ VPWR _03601_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09388_ u_decod.rf_ff_res_data_i\[12\] VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__buf_2
X_08339_ u_rf.reg27_q\[8\] _03365_ _03366_ u_rf.reg19_q\[8\] _03534_ VGND VGND VPWR
+ VPWR _03535_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11350_ _05539_ VGND VGND VPWR VPWR _00887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10301_ u_decod.rf_ff_res_data_i\[18\] VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__buf_2
X_11281_ net531 u_decod.rf_ff_res_data_i\[23\] _05499_ VGND VGND VPWR VPWR _05503_
+ sky130_fd_sc_hd__mux2_1
X_10232_ _04778_ u_rf.reg11_q\[27\] _04922_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__mux2_1
X_10163_ u_rf.reg10_q\[27\] _04484_ _04885_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__mux2_1
X_10094_ _04856_ VGND VGND VPWR VPWR _00314_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_112_clk _00841_ net322 VGND VGND VPWR VPWR u_rf.reg26_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10996_ u_rf.reg22_q\[17\] _04974_ _05344_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12735_ clknet_leaf_136_clk _00772_ net206 VGND VGND VPWR VPWR u_rf.reg24_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12666_ clknet_leaf_93_clk _00703_ net340 VGND VGND VPWR VPWR u_rf.reg21_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12597_ clknet_leaf_46_clk _00634_ net299 VGND VGND VPWR VPWR u_rf.reg19_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11617_ _04766_ u_rf.reg31_q\[21\] _05679_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11548_ _05644_ VGND VGND VPWR VPWR _00980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11479_ _04763_ u_rf.reg29_q\[20\] _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_146_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _02334_ _02908_ _02909_ _02928_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__o31a_2
X_05971_ _01071_ _01247_ _01229_ VGND VGND VPWR VPWR u_decod.dec0.operation_o\[1\]
+ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_29_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08690_ u_rf.reg15_q\[24\] _03301_ _03303_ u_rf.reg24_q\[24\] _03869_ VGND VGND VPWR
+ VPWR _03870_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07641_ _02672_ _02765_ _02766_ _02813_ VGND VGND VPWR VPWR _02863_ sky130_fd_sc_hd__and4_1
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07572_ u_rf.reg9_q\[23\] _02360_ _02386_ u_rf.reg27_q\[23\] _02795_ VGND VGND VPWR
+ VPWR _02796_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06523_ u_rf.reg13_q\[2\] _01598_ _01787_ u_rf.reg18_q\[2\] _01788_ VGND VGND VPWR
+ VPWR _01789_ sky130_fd_sc_hd__a221o_1
X_09311_ _04403_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_146_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09242_ _04355_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06454_ u_rf.reg10_q\[1\] _01656_ _01673_ u_rf.reg2_q\[1\] VGND VGND VPWR VPWR _01722_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09173_ _04297_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06385_ _01513_ _01553_ _01573_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__and3_4
XFILLER_0_113_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08124_ _03241_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08055_ _03257_ VGND VGND VPWR VPWR _03259_ sky130_fd_sc_hd__clkbuf_4
X_07006_ _02189_ _02198_ _02252_ _01505_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_110_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08957_ _04108_ _04111_ VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__xnor2_1
X_07908_ u_rf.reg16_q\[30\] _02307_ _02375_ u_rf.reg11_q\[30\] _03117_ VGND VGND VPWR
+ VPWR _03118_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08888_ _04037_ _04040_ _04045_ _04052_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__a31o_1
X_07839_ _02778_ _02874_ _02964_ _03051_ _01477_ _02685_ VGND VGND VPWR VPWR _03052_
+ sky130_fd_sc_hd__mux4_1
X_10850_ _05274_ VGND VGND VPWR VPWR _00652_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09509_ _04526_ VGND VGND VPWR VPWR _00059_ sky130_fd_sc_hd__clkbuf_1
X_10781_ u_rf.reg19_q\[12\] _04964_ _05235_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__mux2_1
X_12520_ clknet_leaf_59_clk _00557_ net288 VGND VGND VPWR VPWR u_rf.reg17_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12451_ clknet_leaf_108_clk _00488_ net312 VGND VGND VPWR VPWR u_rf.reg15_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11402_ u_rf.reg28_q\[16\] u_decod.rf_ff_res_data_i\[16\] _05560_ VGND VGND VPWR
+ VPWR _05567_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_90 _05319_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_735 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12382_ clknet_leaf_134_clk _00419_ net232 VGND VGND VPWR VPWR u_rf.reg13_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11333_ _05530_ VGND VGND VPWR VPWR _00879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11264_ u_rf.reg26_q\[15\] u_decod.rf_ff_res_data_i\[15\] _05488_ VGND VGND VPWR
+ VPWR _05494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13003_ clknet_leaf_64_clk _01040_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[16\]
+ sky130_fd_sc_hd__dfxtp_2
X_10215_ _04761_ u_rf.reg11_q\[19\] _04911_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__mux2_1
X_11195_ _05457_ VGND VGND VPWR VPWR _00814_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10146_ u_rf.reg10_q\[19\] _04467_ _04874_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10077_ _04847_ VGND VGND VPWR VPWR _00306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10979_ u_rf.reg22_q\[9\] _04957_ _05333_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12718_ clknet_leaf_7_clk _00755_ net218 VGND VGND VPWR VPWR u_rf.reg23_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12649_ clknet_leaf_24_clk _00686_ net266 VGND VGND VPWR VPWR u_rf.reg21_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06170_ u_decod.instr_operation_q\[1\] _01430_ u_decod.instr_unit_q\[1\] _01427_
+ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__o211a_4
XFILLER_0_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09860_ u_rf.reg6_q\[29\] _04488_ _04706_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09791_ u_rf.reg5_q\[29\] _04488_ _04669_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__mux2_1
X_08811_ _03980_ _03982_ _03984_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__or3_1
X_08742_ u_rf.reg18_q\[27\] _03353_ _03355_ u_rf.reg23_q\[27\] _03918_ VGND VGND VPWR
+ VPWR _03919_ sky130_fd_sc_hd__a221o_1
X_05954_ u_decod.dec0.funct3\[0\] VGND VGND VPWR VPWR _01234_ sky130_fd_sc_hd__inv_2
X_08673_ _03844_ _03853_ _03378_ VGND VGND VPWR VPWR _03854_ sky130_fd_sc_hd__o21a_2
X_05885_ u_decod.pc0_q_i\[26\] _01177_ VGND VGND VPWR VPWR _01181_ sky130_fd_sc_hd__or2_1
X_07624_ u_rf.reg22_q\[24\] _01654_ _01668_ u_rf.reg8_q\[24\] VGND VGND VPWR VPWR
+ _02846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07555_ _02734_ _02779_ _02189_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07486_ u_rf.reg29_q\[21\] _01628_ _01639_ u_rf.reg21_q\[21\] _02713_ VGND VGND VPWR
+ VPWR _02714_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06506_ _01713_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__clkbuf_4
X_09225_ _04328_ _04331_ _04336_ _04335_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06437_ _01451_ _01705_ _01500_ VGND VGND VPWR VPWR _01706_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09156_ _04282_ _04283_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06368_ _01637_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__buf_8
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08107_ _03310_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__buf_8
XFILLER_0_114_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09087_ _04223_ _04224_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_110_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_110_clk sky130_fd_sc_hd__clkbuf_16
X_06299_ _01568_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08038_ u_rf.reg28_q\[31\] _03242_ _03243_ u_rf.reg2_q\[31\] VGND VGND VPWR VPWR
+ _03244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_55_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10000_ _04806_ VGND VGND VPWR VPWR _00270_ sky130_fd_sc_hd__clkbuf_1
X_09989_ _04800_ VGND VGND VPWR VPWR _00265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11951_ clknet_leaf_97_clk net490 net332 VGND VGND VPWR VPWR u_decod.pc_q_o\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11882_ clknet_leaf_99_clk u_decod.rs2_data_nxt\[3\] net329 VGND VGND VPWR VPWR u_decod.rs2_data_q\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_10902_ _05302_ VGND VGND VPWR VPWR _00676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10833_ _05265_ VGND VGND VPWR VPWR _00644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10764_ u_rf.reg19_q\[4\] _04947_ _05224_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__mux2_1
X_12503_ clknet_leaf_70_clk _00540_ net352 VGND VGND VPWR VPWR u_rf.reg16_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10695_ _05192_ VGND VGND VPWR VPWR _00579_ sky130_fd_sc_hd__clkbuf_1
X_12434_ clknet_leaf_39_clk _00471_ net277 VGND VGND VPWR VPWR u_rf.reg14_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_770 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_101_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_101_clk sky130_fd_sc_hd__clkbuf_16
X_12365_ clknet_leaf_5_clk _00402_ net215 VGND VGND VPWR VPWR u_rf.reg12_q\[18\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_73_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11316_ _05521_ VGND VGND VPWR VPWR _00871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12296_ clknet_leaf_19_clk _00333_ net282 VGND VGND VPWR VPWR u_rf.reg10_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_11247_ u_rf.reg26_q\[7\] net509 _05477_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
X_11178_ _05448_ VGND VGND VPWR VPWR _00806_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10129_ _04875_ VGND VGND VPWR VPWR _00330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07340_ net199 _02573_ _02489_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09010_ u_decod.rs1_data_q\[28\] u_decod.branch_imm_q_o\[28\] VGND VGND VPWR VPWR
+ _04157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07271_ u_decod.pc_q_o\[17\] _02461_ _02507_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__o21a_1
XFILLER_0_143_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06222_ _01315_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06153_ _01423_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__buf_2
Xhold113 u_exe.pc_data_q\[28\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 u_exe.pc_data_q\[20\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold102 u_decod.flush_v VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 u_decod.rf_ff_res_data_i\[7\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkbuf_2
Xhold157 u_rf.reg26_q\[23\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 u_rf.reg1_q\[20\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__dlygate4sd3_1
X_06084_ _01353_ _01354_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09912_ u_decod.rf_ff_res_data_i\[14\] VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_74_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09843_ _04707_ VGND VGND VPWR VPWR _00212_ sky130_fd_sc_hd__clkbuf_1
X_09774_ _04670_ VGND VGND VPWR VPWR _00180_ sky130_fd_sc_hd__clkbuf_1
X_06986_ _01350_ _01300_ _01304_ _01346_ _02232_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__o41a_1
X_08725_ u_rf.reg31_q\[26\] _03290_ _03292_ u_rf.reg11_q\[26\] _03902_ VGND VGND VPWR
+ VPWR _03903_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05937_ _01071_ _01086_ _01219_ _01094_ VGND VGND VPWR VPWR _01220_ sky130_fd_sc_hd__and4_1
X_08656_ u_rf.reg8_q\[23\] _03407_ _03408_ u_rf.reg29_q\[23\] _03836_ VGND VGND VPWR
+ VPWR _03837_ sky130_fd_sc_hd__a221o_1
X_05868_ u_decod.pc0_q_i\[21\] u_decod.pc0_q_i\[22\] _01162_ VGND VGND VPWR VPWR _01168_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ u_decod.exe_ff_res_data_i\[19\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[19\]
+ _03771_ VGND VGND VPWR VPWR _03772_ sky130_fd_sc_hd__a221o_1
X_07607_ _02681_ _02727_ _02829_ VGND VGND VPWR VPWR _02830_ sky130_fd_sc_hd__o21a_1
X_07538_ u_decod.rf_ff_res_data_i\[22\] _02358_ _02743_ _02744_ _02763_ VGND VGND
+ VPWR VPWR _02764_ sky130_fd_sc_hd__a221o_1
X_05799_ net482 _01105_ _01101_ net92 _01115_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__a221o_1
XFILLER_0_48_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07469_ _01650_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09208_ u_decod.pc_q_o\[22\] u_decod.branch_imm_q_o\[22\] VGND VGND VPWR VPWR _04328_
+ sky130_fd_sc_hd__nand2_1
X_10480_ _04423_ _04568_ _04936_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__or3_4
XFILLER_0_17_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09139_ u_decod.pc_q_o\[12\] u_decod.branch_imm_q_o\[12\] VGND VGND VPWR VPWR _04269_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_20_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12150_ clknet_leaf_48_clk _00187_ net300 VGND VGND VPWR VPWR u_rf.reg5_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11101_ u_rf.reg24_q\[2\] _04943_ _05405_ VGND VGND VPWR VPWR _05408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12081_ clknet_leaf_55_clk _00118_ net294 VGND VGND VPWR VPWR u_rf.reg3_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11032_ _05371_ VGND VGND VPWR VPWR _00737_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ clknet_leaf_70_clk _01020_ net352 VGND VGND VPWR VPWR u_rf.reg31_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11934_ clknet_leaf_79_clk u_decod.rs1_data\[22\] net370 VGND VGND VPWR VPWR u_decod.rs1_data_q\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11865_ clknet_leaf_71_clk _00092_ net358 VGND VGND VPWR VPWR u_rf.reg0_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11796_ clknet_leaf_78_clk net149 net370 VGND VGND VPWR VPWR u_decod.pc0_q_i\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ u_rf.reg19_q\[29\] _04999_ _05246_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10747_ _05219_ VGND VGND VPWR VPWR _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10678_ u_rf.reg17_q\[28\] _04997_ _05174_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12417_ clknet_leaf_118_clk _00454_ net251 VGND VGND VPWR VPWR u_rf.reg14_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12348_ clknet_leaf_127_clk _00385_ net237 VGND VGND VPWR VPWR u_rf.reg12_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12279_ clknet_leaf_50_clk _00316_ net354 VGND VGND VPWR VPWR u_rf.reg9_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06840_ u_decod.rs1_data_q\[9\] _01446_ _01684_ _01753_ VGND VGND VPWR VPWR _02093_
+ sky130_fd_sc_hd__o211a_1
X_06771_ u_rf.reg18_q\[7\] _01590_ _01623_ u_rf.reg28_q\[7\] VGND VGND VPWR VPWR _02027_
+ sky130_fd_sc_hd__a22o_1
X_09490_ _04516_ VGND VGND VPWR VPWR _00050_ sky130_fd_sc_hd__clkbuf_1
X_08510_ u_rf.reg31_q\[16\] _03290_ _03292_ u_rf.reg11_q\[16\] _03697_ VGND VGND VPWR
+ VPWR _03698_ sky130_fd_sc_hd__a221o_1
X_08441_ u_rf.reg16_q\[13\] _03323_ _03313_ u_rf.reg14_q\[13\] _03631_ VGND VGND VPWR
+ VPWR _03632_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08372_ u_rf.reg4_q\[10\] _03265_ _03267_ u_rf.reg17_q\[10\] VGND VGND VPWR VPWR
+ _03566_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07323_ u_rf.reg15_q\[18\] _01601_ _01609_ u_rf.reg12_q\[18\] _02556_ VGND VGND VPWR
+ VPWR _02557_ sky130_fd_sc_hd__a221o_1
X_07254_ _01400_ _01383_ _02443_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__nand3_1
XFILLER_0_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06205_ _01475_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07185_ u_rf.reg3_q\[15\] _02363_ _02364_ u_rf.reg21_q\[15\] _02424_ VGND VGND VPWR
+ VPWR _02425_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_76_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06136_ _01369_ _01399_ _01406_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__or3_2
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06067_ _01307_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _04698_ VGND VGND VPWR VPWR _00204_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ _04661_ VGND VGND VPWR VPWR _00172_ sky130_fd_sc_hd__clkbuf_1
X_06969_ u_rf.reg0_q\[11\] _01663_ _01791_ u_rf.reg10_q\[11\] _02216_ VGND VGND VPWR
+ VPWR _02217_ sky130_fd_sc_hd__a221o_1
X_08708_ u_rf.reg6_q\[25\] _03305_ _03307_ u_rf.reg13_q\[25\] VGND VGND VPWR VPWR
+ _03887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _04623_ VGND VGND VPWR VPWR _00141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08639_ u_rf.reg30_q\[22\] _03200_ _03330_ u_rf.reg28_q\[22\] VGND VGND VPWR VPWR
+ _03821_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11650_ u_decod.branch_imm_q_o\[4\] _01874_ _05696_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _05142_ VGND VGND VPWR VPWR _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11581_ _04730_ u_rf.reg31_q\[4\] _05657_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10532_ _04772_ u_rf.reg15_q\[24\] _05100_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10463_ _05068_ VGND VGND VPWR VPWR _00471_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_118_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10394_ _04770_ u_rf.reg13_q\[23\] _05028_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__mux2_1
X_12202_ clknet_leaf_27_clk _00239_ net266 VGND VGND VPWR VPWR u_rf.reg7_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12133_ clknet_leaf_124_clk _00170_ net231 VGND VGND VPWR VPWR u_rf.reg5_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12064_ clknet_leaf_119_clk _00101_ net247 VGND VGND VPWR VPWR u_rf.reg3_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11015_ u_rf.reg22_q\[26\] _04993_ _05355_ VGND VGND VPWR VPWR _05362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12966_ clknet_leaf_138_clk _01003_ net203 VGND VGND VPWR VPWR u_rf.reg31_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12897_ clknet_leaf_118_clk _00934_ net252 VGND VGND VPWR VPWR u_rf.reg29_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_11917_ clknet_leaf_98_clk u_decod.rs1_data\[5\] net332 VGND VGND VPWR VPWR u_decod.rs1_data_q\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11848_ clknet_leaf_140_clk _00075_ net202 VGND VGND VPWR VPWR u_rf.reg0_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11779_ clknet_leaf_84_clk net162 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08990_ _04132_ _04135_ _04130_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_71_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07941_ u_rf.reg13_q\[31\] _02376_ _01787_ u_rf.reg18_q\[31\] _03148_ VGND VGND VPWR
+ VPWR _03149_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07872_ _01263_ _01266_ _03003_ _01415_ VGND VGND VPWR VPWR _03083_ sky130_fd_sc_hd__a31o_1
X_09611_ _04570_ VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__buf_8
X_06823_ u_rf.reg11_q\[8\] _01582_ _01665_ u_rf.reg8_q\[8\] VGND VGND VPWR VPWR _02077_
+ sky130_fd_sc_hd__a22o_1
X_09542_ u_rf.reg0_q\[10\] _04448_ _04544_ VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__mux2_1
X_06754_ _01335_ _01432_ _02010_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_69_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_102_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ u_rf.reg1_q\[10\] _04448_ _04507_ VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__mux2_1
X_06685_ _01895_ _01899_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__nor2_1
X_08424_ u_rf.reg6_q\[12\] _03305_ _03307_ u_rf.reg13_q\[12\] VGND VGND VPWR VPWR
+ _03616_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08355_ u_rf.reg31_q\[9\] _03290_ _03292_ u_rf.reg11_q\[9\] _03549_ VGND VGND VPWR
+ VPWR _03550_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07306_ _02339_ _02540_ _01458_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08286_ u_rf.reg15_q\[6\] _03300_ _03302_ u_rf.reg24_q\[6\] _03483_ VGND VGND VPWR
+ VPWR _03484_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07237_ u_rf.reg3_q\[16\] _01605_ _01638_ u_rf.reg21_q\[16\] _02474_ VGND VGND VPWR
+ VPWR _02475_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07168_ _01480_ _02351_ _02408_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__a21oi_1
X_06119_ u_decod.rs2_data_q\[16\] _01388_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07099_ net38 _02047_ _02049_ net56 _02051_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout231 net232 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_4
Xfanout220 net255 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net270 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout242 net253 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_2
Xfanout253 net254 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_2
Xfanout275 net276 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_4
Xfanout297 net310 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_2
Xfanout286 net287 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_4
X_09809_ _04689_ VGND VGND VPWR VPWR _00196_ sky130_fd_sc_hd__clkbuf_1
X_12820_ clknet_leaf_22_clk _00857_ net285 VGND VGND VPWR VPWR u_rf.reg26_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12751_ clknet_leaf_35_clk _00788_ net272 VGND VGND VPWR VPWR u_rf.reg24_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11702_ u_decod.branch_imm_q_o\[29\] _03060_ _05717_ VGND VGND VPWR VPWR _05726_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_81_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
X_12682_ clknet_leaf_29_clk _00719_ net259 VGND VGND VPWR VPWR u_rf.reg22_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11633_ _04782_ u_rf.reg31_q\[29\] _05679_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11564_ _05652_ VGND VGND VPWR VPWR _00988_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11495_ _04780_ u_rf.reg29_q\[28\] _05607_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10515_ _04755_ u_rf.reg15_q\[16\] _05089_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_868 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10446_ _05059_ VGND VGND VPWR VPWR _00463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10377_ _04753_ u_rf.reg13_q\[15\] _05017_ VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12116_ clknet_leaf_23_clk _00153_ net267 VGND VGND VPWR VPWR u_rf.reg4_q\[25\] sky130_fd_sc_hd__dfrtp_1
X_12047_ clknet_leaf_73_clk u_decod.exe_ff_res_data_i\[27\] net358 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[27\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12949_ clknet_leaf_54_clk _00986_ net297 VGND VGND VPWR VPWR u_rf.reg30_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06470_ _01234_ _01079_ _01231_ _01083_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__or4_1
XFILLER_0_157_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_191 _03267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_180 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08140_ _03203_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_64_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_846 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08071_ _03274_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__buf_6
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07022_ u_rf.reg11_q\[12\] _01584_ _01598_ u_rf.reg13_q\[12\] _02267_ VGND VGND VPWR
+ VPWR _02268_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08973_ _01367_ u_decod.branch_imm_q_o\[23\] VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__nand2_1
X_07924_ _03130_ _03132_ _01260_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07855_ u_rf.reg7_q\[29\] _01562_ _02363_ u_rf.reg3_q\[29\] VGND VGND VPWR VPWR _03067_
+ sky130_fd_sc_hd__a22o_1
X_07786_ _01264_ _02244_ _03000_ _01820_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__o211a_1
X_06806_ _02059_ _01436_ _02060_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09525_ u_rf.reg0_q\[2\] _04432_ _04533_ VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__mux2_1
X_06737_ u_decod.rs1_data_q\[22\] _01683_ _01292_ u_decod.rs1_data_q\[30\] _01446_
+ _01684_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09456_ u_rf.reg1_q\[2\] _04432_ _04496_ VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__mux2_1
X_06668_ u_rf.reg19_q\[5\] _01593_ _01673_ u_rf.reg2_q\[5\] VGND VGND VPWR VPWR _01928_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08407_ u_rf.reg16_q\[11\] _03450_ _03515_ u_rf.reg5_q\[11\] VGND VGND VPWR VPWR
+ _03600_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06599_ _01860_ _01436_ _01861_ _01435_ _01324_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__a32o_1
X_09387_ _04452_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08338_ u_rf.reg16_q\[8\] _03322_ _03324_ u_rf.reg5_q\[8\] VGND VGND VPWR VPWR _03534_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08269_ u_rf.reg17_q\[5\] _03266_ _03447_ u_rf.reg14_q\[5\] _03467_ VGND VGND VPWR
+ VPWR _03468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11280_ _05502_ VGND VGND VPWR VPWR _00854_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_115_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10300_ _04975_ VGND VGND VPWR VPWR _00401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10231_ _04929_ VGND VGND VPWR VPWR _00378_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_687 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10162_ _04892_ VGND VGND VPWR VPWR _00346_ sky130_fd_sc_hd__clkbuf_1
X_10093_ u_rf.reg9_q\[26\] _04482_ _04849_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12803_ clknet_leaf_106_clk _00840_ net320 VGND VGND VPWR VPWR u_rf.reg26_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_54_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12734_ clknet_leaf_134_clk _00771_ net209 VGND VGND VPWR VPWR u_rf.reg24_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ _05351_ VGND VGND VPWR VPWR _00720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12665_ clknet_leaf_64_clk _00702_ net341 VGND VGND VPWR VPWR u_rf.reg21_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11616_ _05680_ VGND VGND VPWR VPWR _01012_ sky130_fd_sc_hd__clkbuf_1
X_12596_ clknet_leaf_32_clk _00633_ net263 VGND VGND VPWR VPWR u_rf.reg19_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_13_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11547_ _04763_ u_rf.reg30_q\[20\] _05643_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11478_ _05584_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__buf_6
X_10429_ _05050_ VGND VGND VPWR VPWR _00455_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05970_ _01090_ _01221_ _01246_ _01084_ _01244_ VGND VGND VPWR VPWR _01247_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_146_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07640_ _01528_ _02840_ _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__o21a_1
X_07571_ u_rf.reg12_q\[23\] _01609_ _01674_ u_rf.reg2_q\[23\] VGND VGND VPWR VPWR
+ _02795_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_45_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06522_ u_rf.reg30_q\[2\] _01580_ _01625_ u_rf.reg28_q\[2\] VGND VGND VPWR VPWR _01788_
+ sky130_fd_sc_hd__a22o_1
X_09310_ _04397_ u_decod.rs2_data_q\[17\] _04398_ VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_66_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09241_ u_decod.pc_q_o\[27\] u_decod.branch_imm_q_o\[27\] VGND VGND VPWR VPWR _04356_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_806 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06453_ u_rf.reg1_q\[1\] _01586_ _01615_ u_rf.reg31_q\[1\] _01720_ VGND VGND VPWR
+ VPWR _01721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09172_ _04283_ _04287_ _04291_ _04290_ VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06384_ _01653_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__buf_6
XFILLER_0_43_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08123_ u_rf.reg27_q\[0\] _03319_ _03321_ u_rf.reg19_q\[0\] _03326_ VGND VGND VPWR
+ VPWR _03327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08054_ _03258_ VGND VGND VPWR VPWR u_decod.rs1_data_nxt\[32\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07005_ _01479_ _02251_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08956_ _04096_ _04099_ _04103_ _04110_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__o31a_1
XPHY_EDGE_ROW_102_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07907_ u_rf.reg15_q\[30\] _02371_ _01654_ u_rf.reg22_q\[30\] VGND VGND VPWR VPWR
+ _03117_ sky130_fd_sc_hd__a22o_1
X_08887_ u_decod.rs1_data_q\[8\] u_decod.branch_imm_q_o\[8\] _04051_ _04044_ VGND
+ VGND VPWR VPWR _04052_ sky130_fd_sc_hd__a31o_1
X_07838_ u_decod.rs1_data_q\[29\] _01358_ u_decod.rs1_data_q\[13\] u_decod.rs1_data_q\[5\]
+ _01469_ _01466_ VGND VGND VPWR VPWR _03051_ sky130_fd_sc_hd__mux4_1
X_09508_ u_rf.reg1_q\[27\] _04484_ _04518_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__mux2_1
X_07769_ u_rf.reg7_q\[27\] _01562_ _02363_ u_rf.reg3_q\[27\] VGND VGND VPWR VPWR _02985_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_36_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10780_ _05237_ VGND VGND VPWR VPWR _00619_ sky130_fd_sc_hd__clkbuf_1
X_09439_ _04487_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12450_ clknet_leaf_130_clk _00487_ net229 VGND VGND VPWR VPWR u_rf.reg15_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11401_ _05566_ VGND VGND VPWR VPWR _00911_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_91 _05427_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_80 _04838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12381_ clknet_leaf_15_clk _00418_ net245 VGND VGND VPWR VPWR u_rf.reg13_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11332_ _04753_ u_rf.reg27_q\[15\] _05524_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11263_ _05493_ VGND VGND VPWR VPWR _00846_ sky130_fd_sc_hd__clkbuf_1
X_11194_ u_rf.reg25_q\[14\] _04968_ _05452_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__mux2_1
X_13002_ clknet_leaf_92_clk _01039_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[15\]
+ sky130_fd_sc_hd__dfxtp_2
X_10214_ _04920_ VGND VGND VPWR VPWR _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10145_ _04883_ VGND VGND VPWR VPWR _00338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_392 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ u_rf.reg9_q\[18\] _04465_ _04838_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_18_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10978_ _05342_ VGND VGND VPWR VPWR _00712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12717_ clknet_leaf_5_clk _00754_ net217 VGND VGND VPWR VPWR u_rf.reg23_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12648_ clknet_leaf_17_clk _00685_ net289 VGND VGND VPWR VPWR u_rf.reg21_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12579_ clknet_leaf_109_clk _00616_ net313 VGND VGND VPWR VPWR u_rf.reg19_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_635 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08810_ u_rf.reg8_q\[30\] _03270_ _03272_ u_rf.reg29_q\[30\] _03983_ VGND VGND VPWR
+ VPWR _03984_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09790_ _04678_ VGND VGND VPWR VPWR _00188_ sky130_fd_sc_hd__clkbuf_1
X_08741_ u_rf.reg4_q\[27\] _03265_ _03267_ u_rf.reg17_q\[27\] VGND VGND VPWR VPWR
+ _03918_ sky130_fd_sc_hd__a22o_1
X_05953_ _01231_ _01085_ _01209_ _01232_ VGND VGND VPWR VPWR _01233_ sky130_fd_sc_hd__or4_1
X_08672_ _03846_ _03848_ _03850_ _03852_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__or4_1
X_05884_ u_decod.pc0_q_i\[26\] _01177_ VGND VGND VPWR VPWR _01180_ sky130_fd_sc_hd__and2_4
X_07623_ u_rf.reg6_q\[24\] _01557_ _02376_ u_rf.reg13_q\[24\] _02844_ VGND VGND VPWR
+ VPWR _02845_ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07554_ _02498_ _02584_ _02684_ _02778_ _01476_ _02685_ VGND VGND VPWR VPWR _02779_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07485_ u_rf.reg1_q\[21\] _01587_ _01659_ u_rf.reg14_q\[21\] VGND VGND VPWR VPWR
+ _02713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06505_ _01746_ _01751_ _01760_ _01771_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[2\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09224_ _04340_ _04341_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06436_ _01455_ _01704_ _01497_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__o21a_1
XFILLER_0_16_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09155_ u_decod.pc_q_o\[14\] u_decod.branch_imm_q_o\[14\] VGND VGND VPWR VPWR _04283_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06367_ _01572_ _01566_ _01551_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__and3_2
X_08106_ _03231_ VGND VGND VPWR VPWR _03310_ sky130_fd_sc_hd__buf_8
X_09086_ _04210_ _04215_ _04214_ _04216_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06298_ _01567_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08037_ _03170_ _03173_ _03199_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09988_ u_rf.reg8_q\[9\] _04446_ _04790_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__mux2_1
X_08939_ _04094_ _04095_ VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11950_ clknet_leaf_117_clk u_decod.dec0.rd_o\[4\] net325 VGND VGND VPWR VPWR u_decod.exe_ff_rd_adr_q_i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ u_rf.reg21_q\[4\] _04947_ _05297_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[2\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10832_ u_rf.reg20_q\[4\] _04947_ _05260_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10763_ _05228_ VGND VGND VPWR VPWR _00611_ sky130_fd_sc_hd__clkbuf_1
X_12502_ clknet_leaf_47_clk _00539_ net300 VGND VGND VPWR VPWR u_rf.reg16_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10694_ u_rf.reg18_q\[3\] _04945_ _05188_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__mux2_1
X_12433_ clknet_leaf_54_clk _00470_ net302 VGND VGND VPWR VPWR u_rf.reg14_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12364_ clknet_leaf_20_clk _00401_ net280 VGND VGND VPWR VPWR u_rf.reg12_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11315_ _04736_ u_rf.reg27_q\[7\] _05513_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_432 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12295_ clknet_leaf_4_clk _00332_ net212 VGND VGND VPWR VPWR u_rf.reg10_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11246_ _05484_ VGND VGND VPWR VPWR _00838_ sky130_fd_sc_hd__clkbuf_1
X_11177_ u_rf.reg25_q\[6\] _04951_ _05441_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__mux2_1
X_10128_ u_rf.reg10_q\[10\] _04448_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10059_ _04826_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__buf_8
XFILLER_0_89_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07270_ _02334_ _02506_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06221_ net33 _01487_ _01488_ net40 _01491_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_413 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06152_ _01422_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_4
Xhold125 u_exe.pc_data_q\[25\] VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 u_decod.rf_ff_res_data_i\[24\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold114 u_exe.pc_data_q\[12\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__dlygate4sd3_1
X_06083_ u_decod.rs2_data_q\[14\] _01292_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold136 u_exe.pc_data_q\[30\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09911_ _04750_ VGND VGND VPWR VPWR _00237_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_7_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold147 u_rf.reg19_q\[16\] VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09842_ u_rf.reg6_q\[20\] _04469_ _04706_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__mux2_1
X_09773_ u_rf.reg5_q\[20\] _04469_ _04669_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__mux2_1
X_08724_ u_rf.reg9_q\[26\] _03294_ _03296_ u_rf.reg20_q\[26\] VGND VGND VPWR VPWR
+ _03902_ sky130_fd_sc_hd__a22o_1
X_06985_ _02231_ _01436_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__and2_1
X_05936_ _01080_ u_decod.dec0.funct7\[6\] _01082_ VGND VGND VPWR VPWR _01219_ sky130_fd_sc_hd__nor3_1
X_08655_ u_rf.reg22_q\[23\] _03274_ _03410_ u_rf.reg3_q\[23\] VGND VGND VPWR VPWR
+ _03836_ sky130_fd_sc_hd__a22o_1
X_05867_ _01099_ _01165_ _01166_ _01167_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__a31o_1
XFILLER_0_96_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03754_ _03763_ _03770_ _03253_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__o31a_2
X_07606_ _02681_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__nand2_1
X_07537_ _02753_ _02762_ _02359_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__o21a_1
X_05798_ _01113_ _01106_ _01114_ VGND VGND VPWR VPWR _01115_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07468_ u_decod.dec0.instr_i\[21\] _01206_ _02645_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09207_ _04116_ _04274_ _04275_ _04327_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[21\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_107_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07399_ _02449_ _02629_ _01905_ VGND VGND VPWR VPWR _02630_ sky130_fd_sc_hd__mux2_1
X_06419_ _01315_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09138_ u_decod.pc_q_o\[12\] u_decod.branch_imm_q_o\[12\] VGND VGND VPWR VPWR _04268_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_17_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09069_ _04198_ _04202_ _04203_ VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11100_ _05407_ VGND VGND VPWR VPWR _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12080_ clknet_leaf_36_clk _00117_ net271 VGND VGND VPWR VPWR u_rf.reg3_q\[21\] sky130_fd_sc_hd__dfrtp_1
X_11031_ _04724_ u_rf.reg23_q\[1\] _05369_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ clknet_leaf_49_clk _01019_ net309 VGND VGND VPWR VPWR u_rf.reg31_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_11933_ clknet_leaf_79_clk u_decod.rs1_data\[21\] net371 VGND VGND VPWR VPWR u_decod.rs1_data_q\[21\]
+ sky130_fd_sc_hd__dfrtp_2
X_11864_ clknet_leaf_51_clk _00091_ net307 VGND VGND VPWR VPWR u_rf.reg0_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10815_ _05255_ VGND VGND VPWR VPWR _00636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_830 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ clknet_leaf_78_clk net148 net370 VGND VGND VPWR VPWR u_decod.pc0_q_i\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10746_ u_rf.reg18_q\[28\] _04997_ _05210_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10677_ _05182_ VGND VGND VPWR VPWR _00571_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12416_ clknet_leaf_120_clk _00453_ net248 VGND VGND VPWR VPWR u_rf.reg14_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12347_ clknet_leaf_12_clk _00384_ net243 VGND VGND VPWR VPWR u_rf.reg12_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12278_ clknet_leaf_51_clk _00315_ net308 VGND VGND VPWR VPWR u_rf.reg9_q\[27\] sky130_fd_sc_hd__dfrtp_1
X_11229_ u_rf.reg25_q\[31\] _05003_ _05440_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06770_ u_rf.reg19_q\[7\] _01594_ _01627_ u_rf.reg29_q\[7\] _02025_ VGND VGND VPWR
+ VPWR _02026_ sky130_fd_sc_hd__a221o_1
X_08440_ u_rf.reg31_q\[13\] _03289_ _03285_ u_rf.reg21_q\[13\] VGND VGND VPWR VPWR
+ _03631_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08371_ _03257_ VGND VGND VPWR VPWR _03565_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07322_ u_rf.reg25_q\[18\] _01576_ _01625_ u_rf.reg28_q\[18\] VGND VGND VPWR VPWR
+ _02556_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07253_ _01400_ _02443_ _01383_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_104_719 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07184_ u_rf.reg5_q\[15\] _01569_ _01556_ u_rf.reg6_q\[15\] VGND VGND VPWR VPWR _02424_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06204_ _01474_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__buf_4
X_06135_ _01375_ _01405_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06066_ _01306_ _01305_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__nor2_1
X_09825_ u_rf.reg6_q\[12\] _04453_ _04695_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ u_rf.reg5_q\[12\] _04453_ _04658_ VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__mux2_1
X_06968_ u_rf.reg29_q\[11\] _01627_ _01658_ u_rf.reg14_q\[11\] VGND VGND VPWR VPWR
+ _02216_ sky130_fd_sc_hd__a22o_1
X_08707_ u_rf.reg7_q\[25\] _03369_ _03370_ u_rf.reg25_q\[25\] _03885_ VGND VGND VPWR
+ VPWR _03886_ sky130_fd_sc_hd__a221o_1
X_09687_ u_rf.reg4_q\[13\] _04455_ _04619_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__mux2_1
X_05919_ _01079_ _01082_ VGND VGND VPWR VPWR _01209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ u_rf.reg22_q\[22\] _03275_ _03270_ u_rf.reg8_q\[22\] _03819_ VGND VGND VPWR
+ VPWR _03820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ u_decod.pc_q_o\[9\] u_decod.pc_q_o\[10\] _02054_ VGND VGND VPWR VPWR _02150_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08569_ u_rf.reg0_q\[19\] _03176_ _03329_ u_rf.reg12_q\[19\] _03753_ VGND VGND VPWR
+ VPWR _03754_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_25_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10600_ u_rf.reg16_q\[23\] _04987_ _05138_ VGND VGND VPWR VPWR _05142_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11580_ _05661_ VGND VGND VPWR VPWR _00995_ sky130_fd_sc_hd__clkbuf_1
X_10531_ _05104_ VGND VGND VPWR VPWR _00503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_360 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10462_ _04770_ u_rf.reg14_q\[23\] _05064_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ clknet_leaf_19_clk _00238_ net281 VGND VGND VPWR VPWR u_rf.reg7_q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_875 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10393_ _05031_ VGND VGND VPWR VPWR _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12132_ clknet_leaf_111_clk _00169_ net316 VGND VGND VPWR VPWR u_rf.reg5_q\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12063_ clknet_leaf_131_clk _00100_ net227 VGND VGND VPWR VPWR u_rf.reg3_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11014_ _05361_ VGND VGND VPWR VPWR _00729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12965_ clknet_leaf_126_clk _01002_ net240 VGND VGND VPWR VPWR u_rf.reg31_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11916_ clknet_leaf_102_clk u_decod.rs1_data\[4\] net337 VGND VGND VPWR VPWR u_decod.rs1_data_q\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12896_ clknet_leaf_120_clk _00933_ net324 VGND VGND VPWR VPWR u_rf.reg29_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11847_ clknet_leaf_121_clk _00074_ net247 VGND VGND VPWR VPWR u_rf.reg0_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11778_ clknet_leaf_87_clk net161 net362 VGND VGND VPWR VPWR u_decod.pc0_q_i\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10729_ _05187_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07940_ u_rf.reg27_q\[31\] _02386_ _01776_ u_rf.reg2_q\[31\] VGND VGND VPWR VPWR
+ _03148_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07871_ _03081_ _03082_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[29\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09610_ _04581_ VGND VGND VPWR VPWR _00105_ sky130_fd_sc_hd__clkbuf_1
X_06822_ u_rf.reg0_q\[8\] _01516_ _01599_ u_rf.reg15_q\[8\] _02075_ VGND VGND VPWR
+ VPWR _02076_ sky130_fd_sc_hd__a221o_1
X_09541_ _04532_ VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__buf_8
X_06753_ _01326_ _01429_ _01435_ _01327_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09472_ _04495_ VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_69_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06684_ _01713_ u_decod.exe_ff_res_data_i\[5\] _01943_ VGND VGND VPWR VPWR _01944_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08423_ _03608_ _03610_ _03612_ _03614_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08354_ u_rf.reg9_q\[9\] _03294_ _03296_ u_rf.reg20_q\[9\] VGND VGND VPWR VPWR _03549_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07305_ _01384_ _01302_ u_decod.rs1_data_q\[2\] _01747_ _01455_ _01447_ VGND VGND
+ VPWR VPWR _02540_ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08285_ u_rf.reg6_q\[6\] _03304_ _03306_ u_rf.reg13_q\[6\] VGND VGND VPWR VPWR _03483_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07236_ u_rf.reg5_q\[16\] _01568_ _01555_ u_rf.reg6_q\[16\] VGND VGND VPWR VPWR _02474_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07167_ _01480_ _02407_ _01442_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06118_ u_decod.rs2_data_q\[16\] _01388_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07098_ _02292_ _02249_ _02295_ _02340_ _01480_ _01477_ VGND VGND VPWR VPWR _02341_
+ sky130_fd_sc_hd__mux4_2
X_06049_ u_decod.rs1_data_q\[3\] u_decod.rs2_data_q\[3\] VGND VGND VPWR VPWR _01320_
+ sky130_fd_sc_hd__nand2_1
Xfanout221 net223 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_4
Xfanout210 net255 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__buf_2
Xfanout232 net233 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout265 net266 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net253 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_4
Xfanout254 net255 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_2
Xfanout298 net301 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_4
Xfanout276 net311 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__buf_2
Xfanout287 net310 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_89_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09808_ u_rf.reg6_q\[4\] _04436_ _04684_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09739_ u_rf.reg5_q\[4\] _04436_ _04647_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12750_ clknet_leaf_29_clk _00787_ net256 VGND VGND VPWR VPWR u_rf.reg24_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11701_ _05725_ VGND VGND VPWR VPWR _01052_ sky130_fd_sc_hd__clkbuf_1
X_12681_ clknet_leaf_24_clk _00718_ net267 VGND VGND VPWR VPWR u_rf.reg22_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11632_ _05688_ VGND VGND VPWR VPWR _01020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11563_ _04780_ u_rf.reg30_q\[28\] _05643_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11494_ _05615_ VGND VGND VPWR VPWR _00955_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ _05095_ VGND VGND VPWR VPWR _00495_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10445_ _04753_ u_rf.reg14_q\[15\] _05053_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12115_ clknet_leaf_53_clk _00152_ net304 VGND VGND VPWR VPWR u_rf.reg4_q\[24\] sky130_fd_sc_hd__dfrtp_1
X_10376_ _05022_ VGND VGND VPWR VPWR _00430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12046_ clknet_leaf_74_clk u_decod.exe_ff_res_data_i\[26\] net356 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[26\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_148_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_148_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_23_clk _00985_ net284 VGND VGND VPWR VPWR u_rf.reg30_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12879_ clknet_leaf_44_clk _00916_ net295 VGND VGND VPWR VPWR u_rf.reg28_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_170 u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_192 _03267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_157_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08070_ _03218_ VGND VGND VPWR VPWR _03274_ sky130_fd_sc_hd__buf_8
XFILLER_0_55_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07021_ u_rf.reg30_q\[12\] _01579_ _01591_ u_rf.reg18_q\[12\] VGND VGND VPWR VPWR
+ _02267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08972_ _01367_ u_decod.branch_imm_q_o\[23\] VGND VGND VPWR VPWR _04124_ sky130_fd_sc_hd__or2_1
X_07923_ _01269_ _03131_ _02781_ _01268_ VGND VGND VPWR VPWR _03132_ sky130_fd_sc_hd__a2bb2o_1
X_07854_ u_rf.reg25_q\[29\] _01783_ _02652_ u_rf.reg23_q\[29\] _03065_ VGND VGND VPWR
+ VPWR _03066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06805_ _01340_ _01332_ _01336_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__or3_1
X_07785_ _02781_ _01264_ VGND VGND VPWR VPWR _03000_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09524_ _04535_ VGND VGND VPWR VPWR _00065_ sky130_fd_sc_hd__clkbuf_1
X_06736_ _01327_ _01992_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06667_ u_rf.reg25_q\[5\] _01575_ _01670_ u_rf.reg27_q\[5\] _01926_ VGND VGND VPWR
+ VPWR _01927_ sky130_fd_sc_hd__a221o_1
X_09455_ _04498_ VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08406_ u_rf.reg7_q\[11\] _03428_ _03429_ u_rf.reg25_q\[11\] _03598_ VGND VGND VPWR
+ VPWR _03599_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06598_ _01321_ _01324_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__or2_1
X_09386_ u_rf.reg2_q\[11\] _04451_ _04449_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08337_ u_rf.reg0_q\[8\] _03175_ _03421_ u_rf.reg12_q\[8\] _03532_ VGND VGND VPWR
+ VPWR _03533_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08268_ u_rf.reg28_q\[5\] _03330_ _03332_ u_rf.reg2_q\[5\] VGND VGND VPWR VPWR _03467_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07219_ _01688_ _02456_ _02457_ _01478_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__a211o_1
X_10230_ _04776_ u_rf.reg11_q\[26\] _04922_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__mux2_1
X_08199_ u_rf.reg18_q\[2\] _03352_ _03354_ u_rf.reg23_q\[2\] _03400_ VGND VGND VPWR
+ VPWR _03401_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10161_ u_rf.reg10_q\[26\] _04482_ _04885_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__mux2_1
X_10092_ _04855_ VGND VGND VPWR VPWR _00313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12802_ clknet_leaf_129_clk _00839_ net235 VGND VGND VPWR VPWR u_rf.reg26_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10994_ u_rf.reg22_q\[16\] _04972_ _05344_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_815 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12733_ clknet_leaf_19_clk _00770_ net281 VGND VGND VPWR VPWR u_rf.reg24_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12664_ clknet_leaf_64_clk _00701_ net342 VGND VGND VPWR VPWR u_rf.reg21_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12595_ clknet_leaf_69_clk _00632_ net350 VGND VGND VPWR VPWR u_rf.reg19_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11615_ _04763_ u_rf.reg31_q\[20\] _05679_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11546_ _05620_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11477_ _05606_ VGND VGND VPWR VPWR _00947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10428_ _04736_ u_rf.reg14_q\[7\] _05042_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10359_ _05013_ VGND VGND VPWR VPWR _00422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12029_ clknet_leaf_113_clk u_decod.exe_ff_res_data_i\[9\] net322 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_23 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07570_ u_rf.reg31_q\[23\] _01777_ _02697_ u_rf.reg4_q\[23\] _02793_ VGND VGND VPWR
+ VPWR _02794_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06521_ _01592_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09240_ u_decod.pc_q_o\[27\] u_decod.branch_imm_q_o\[27\] VGND VGND VPWR VPWR _04355_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06452_ u_rf.reg28_q\[1\] _01624_ _01644_ u_rf.reg20_q\[1\] VGND VGND VPWR VPWR _01720_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09171_ _04295_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06383_ _01652_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__buf_6
XFILLER_0_44_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08122_ u_rf.reg16_q\[0\] _03323_ _03325_ u_rf.reg5_q\[0\] VGND VGND VPWR VPWR _03326_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08053_ u_decod.dec0.unsign_extension u_decod.rs1_data\[31\] VGND VGND VPWR VPWR
+ _03258_ sky130_fd_sc_hd__and2b_1
XFILLER_0_114_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07004_ _02144_ _02250_ _01474_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08955_ _01376_ u_decod.branch_imm_q_o\[19\] _04109_ VGND VGND VPWR VPWR _04110_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_110_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07906_ u_rf.reg6_q\[30\] _01557_ _02697_ u_rf.reg4_q\[30\] _03115_ VGND VGND VPWR
+ VPWR _03116_ sky130_fd_sc_hd__a221o_1
X_08886_ u_decod.rs1_data_q\[9\] u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _04051_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07837_ _02619_ net54 _02618_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__a21bo_1
X_07768_ u_rf.reg5_q\[27\] _02664_ _02665_ u_rf.reg19_q\[27\] _02983_ VGND VGND VPWR
+ VPWR _02984_ sky130_fd_sc_hd__a221o_1
X_09507_ _04525_ VGND VGND VPWR VPWR _00058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06719_ _01970_ _01972_ _01974_ _01976_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07699_ _02732_ _02917_ _02685_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09438_ u_rf.reg2_q\[28\] _04486_ _04470_ VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09369_ u_decod.rf_ff_res_data_i\[6\] VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11400_ u_rf.reg28_q\[15\] u_decod.rf_ff_res_data_i\[15\] _05560_ VGND VGND VPWR
+ VPWR _05566_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12380_ clknet_leaf_126_clk _00417_ net240 VGND VGND VPWR VPWR u_rf.reg13_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_70 _04518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11331_ _05529_ VGND VGND VPWR VPWR _00878_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_92 _05441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _04838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11262_ u_rf.reg26_q\[14\] u_decod.rf_ff_res_data_i\[14\] _05488_ VGND VGND VPWR
+ VPWR _05493_ sky130_fd_sc_hd__mux2_1
X_13001_ clknet_leaf_92_clk _01038_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[14\]
+ sky130_fd_sc_hd__dfxtp_2
X_11193_ _05456_ VGND VGND VPWR VPWR _00813_ sky130_fd_sc_hd__clkbuf_1
X_10213_ _04759_ u_rf.reg11_q\[18\] _04911_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10144_ u_rf.reg10_q\[18\] _04465_ _04874_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ _04846_ VGND VGND VPWR VPWR _00305_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10977_ u_rf.reg22_q\[8\] _04955_ _05333_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12716_ clknet_leaf_10_clk _00753_ net224 VGND VGND VPWR VPWR u_rf.reg23_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ clknet_leaf_3_clk _00684_ net211 VGND VGND VPWR VPWR u_rf.reg21_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12578_ clknet_leaf_132_clk _00615_ net230 VGND VGND VPWR VPWR u_rf.reg19_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11529_ _05634_ VGND VGND VPWR VPWR _00971_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08740_ u_rf.reg8_q\[27\] _03407_ _03408_ u_rf.reg29_q\[27\] _03916_ VGND VGND VPWR
+ VPWR _03917_ sky130_fd_sc_hd__a221o_1
X_05952_ _01080_ u_decod.dec0.funct3\[0\] u_decod.dec0.funct7\[6\] VGND VGND VPWR
+ VPWR _01232_ sky130_fd_sc_hd__or3_1
X_08671_ u_rf.reg28_q\[23\] _03331_ _03333_ u_rf.reg2_q\[23\] _03851_ VGND VGND VPWR
+ VPWR _03852_ sky130_fd_sc_hd__a221o_1
X_05883_ net499 _01142_ _01132_ net82 _01179_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__a221o_1
XFILLER_0_84_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07622_ u_rf.reg30_q\[24\] _01581_ _01636_ u_rf.reg9_q\[24\] VGND VGND VPWR VPWR
+ _02844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_494 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07553_ _01367_ _01289_ u_decod.rs1_data_q\[7\] _01747_ _01468_ _01466_ VGND VGND
+ VPWR VPWR _02778_ sky130_fd_sc_hd__mux4_1
X_07484_ u_rf.reg25_q\[21\] _01576_ _01622_ u_rf.reg24_q\[21\] _02711_ VGND VGND VPWR
+ VPWR _02712_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06504_ _01059_ _01762_ _01768_ _01770_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__a211o_1
X_09223_ u_decod.pc_q_o\[24\] u_decod.branch_imm_q_o\[24\] VGND VGND VPWR VPWR _04341_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_124_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06435_ net409 _01702_ _01703_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__o21a_1
X_09154_ u_decod.pc_q_o\[14\] u_decod.branch_imm_q_o\[14\] VGND VGND VPWR VPWR _04282_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_745 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08105_ u_rf.reg15_q\[0\] _03301_ _03303_ u_rf.reg24_q\[0\] _03308_ VGND VGND VPWR
+ VPWR _03309_ sky130_fd_sc_hd__a221o_1
X_06366_ _01635_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09085_ _04221_ _04222_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06297_ _01513_ _01566_ _01551_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__and3_2
XFILLER_0_141_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08036_ u_decod.dec0.instr_i\[19\] _03172_ _03198_ VGND VGND VPWR VPWR _03242_ sky130_fd_sc_hd__and3_2
Xinput90 reset_adr_i[3] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XFILLER_0_31_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09987_ _04799_ VGND VGND VPWR VPWR _00264_ sky130_fd_sc_hd__clkbuf_1
X_08938_ _01384_ u_decod.branch_imm_q_o\[18\] VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__nand2_1
X_08869_ u_decod.rs1_data_q\[8\] u_decod.branch_imm_q_o\[8\] VGND VGND VPWR VPWR _04036_
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_4_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _05301_ VGND VGND VPWR VPWR _00675_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_123_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11880_ clknet_leaf_113_clk u_decod.rs2_data_nxt\[1\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_123_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10831_ _05264_ VGND VGND VPWR VPWR _00643_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10762_ u_rf.reg19_q\[3\] _04945_ _05224_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12501_ clknet_leaf_46_clk _00538_ net298 VGND VGND VPWR VPWR u_rf.reg16_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12432_ clknet_leaf_36_clk _00469_ net273 VGND VGND VPWR VPWR u_rf.reg14_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10693_ _05191_ VGND VGND VPWR VPWR _00578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12363_ clknet_leaf_1_clk _00400_ net208 VGND VGND VPWR VPWR u_rf.reg12_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_11314_ _05520_ VGND VGND VPWR VPWR _00870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12294_ clknet_leaf_140_clk _00331_ net202 VGND VGND VPWR VPWR u_rf.reg10_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11245_ u_rf.reg26_q\[6\] u_decod.rf_ff_res_data_i\[6\] _05477_ VGND VGND VPWR VPWR
+ _05484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11176_ _05447_ VGND VGND VPWR VPWR _00805_ sky130_fd_sc_hd__clkbuf_1
X_10127_ _04862_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__buf_8
XFILLER_0_145_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10058_ _04837_ VGND VGND VPWR VPWR _00297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_121_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06220_ net63 _01489_ _01490_ net49 VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_130_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06151_ u_decod.rs2_data_q\[0\] VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 u_exe.pc_data_q\[19\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 u_exe.pc_data_q\[31\] VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold104 u_exe.pc_data_q\[7\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06082_ u_decod.rs2_data_q\[14\] _01292_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__and2_1
X_09910_ _04749_ u_rf.reg7_q\[13\] _04743_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__mux2_1
Xhold137 u_decod.dec0.instr_i\[8\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold148 u_rf.reg6_q\[1\] VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09841_ _04683_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09772_ _04646_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__buf_6
X_06984_ _01300_ _01304_ _01346_ _01350_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__o31ai_1
X_08723_ u_rf.reg30_q\[26\] _03280_ _03282_ u_rf.reg10_q\[26\] _03900_ VGND VGND VPWR
+ VPWR _03901_ sky130_fd_sc_hd__a221o_1
X_05935_ _01068_ _01201_ _01070_ VGND VGND VPWR VPWR u_decod.dec0.is_branch sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05866_ net517 _01118_ _01119_ net78 VGND VGND VPWR VPWR _01167_ sky130_fd_sc_hd__a22o_1
X_08654_ net438 _03773_ _03835_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[22\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05797_ u_decod.pc0_q_i\[5\] _01110_ VGND VGND VPWR VPWR _01114_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08585_ _03765_ _03767_ _03769_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__or3_1
X_07605_ _02623_ _02827_ _01472_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__mux2_1
X_07536_ _02755_ _02757_ _02759_ _02761_ VGND VGND VPWR VPWR _02762_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09206_ _04325_ _04326_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__xnor2_1
X_07467_ _02695_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[21\] sky130_fd_sc_hd__inv_2
XFILLER_0_151_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07398_ _01363_ _01297_ u_decod.rs1_data_q\[4\] _01747_ _01460_ _01461_ VGND VGND
+ VPWR VPWR _02629_ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06418_ _01471_ _01686_ _01464_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09137_ _04059_ _04207_ _04208_ _04267_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[11\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06349_ _01571_ _01589_ _01603_ _01618_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09068_ _04196_ VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__buf_2
X_08019_ _03188_ _03173_ _03204_ VGND VGND VPWR VPWR _03225_ sky130_fd_sc_hd__and3_4
XFILLER_0_130_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11030_ _05370_ VGND VGND VPWR VPWR _00736_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_125_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12981_ clknet_leaf_45_clk _01018_ net298 VGND VGND VPWR VPWR u_rf.reg31_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_11932_ clknet_leaf_80_clk u_decod.rs1_data\[20\] net371 VGND VGND VPWR VPWR u_decod.rs1_data_q\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11863_ clknet_leaf_44_clk _00090_ net296 VGND VGND VPWR VPWR u_rf.reg0_q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10814_ u_rf.reg19_q\[28\] _04997_ _05246_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11794_ clknet_leaf_78_clk net147 net370 VGND VGND VPWR VPWR u_decod.pc0_q_i\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10745_ _05218_ VGND VGND VPWR VPWR _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10676_ u_rf.reg17_q\[27\] _04995_ _05174_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12415_ clknet_leaf_132_clk _00452_ net227 VGND VGND VPWR VPWR u_rf.reg14_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_388 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12346_ clknet_leaf_61_clk _00383_ net341 VGND VGND VPWR VPWR u_rf.reg11_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12277_ clknet_leaf_44_clk _00314_ net294 VGND VGND VPWR VPWR u_rf.reg9_q\[26\] sky130_fd_sc_hd__dfrtp_1
X_11228_ _05474_ VGND VGND VPWR VPWR _00830_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11159_ u_rf.reg24_q\[30\] _05001_ _05404_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08370_ net465 _03259_ _03564_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[9\]
+ sky130_fd_sc_hd__a22o_1
X_07321_ u_rf.reg19_q\[18\] _01595_ _01650_ u_rf.reg4_q\[18\] _02554_ VGND VGND VPWR
+ VPWR _02555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07252_ _02486_ _02489_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[16\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07183_ u_rf.reg31_q\[15\] _01616_ _02367_ u_rf.reg14_q\[15\] _02422_ VGND VGND VPWR
+ VPWR _02423_ sky130_fd_sc_hd__a221o_1
X_06203_ _01315_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06134_ _01377_ _01404_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__nand2_2
XFILLER_0_53_191 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06065_ _01326_ _01329_ _01334_ _01335_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__o31a_1
XFILLER_0_1_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09824_ _04697_ VGND VGND VPWR VPWR _00203_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _04660_ VGND VGND VPWR VPWR _00171_ sky130_fd_sc_hd__clkbuf_1
X_06967_ u_rf.reg25_q\[11\] _01576_ _01580_ u_rf.reg30_q\[11\] _02214_ VGND VGND VPWR
+ VPWR _02215_ sky130_fd_sc_hd__a221o_1
X_08706_ u_rf.reg1_q\[25\] _03310_ _03312_ u_rf.reg14_q\[25\] VGND VGND VPWR VPWR
+ _03885_ sky130_fd_sc_hd__a22o_1
X_09686_ _04622_ VGND VGND VPWR VPWR _00140_ sky130_fd_sc_hd__clkbuf_1
X_06898_ u_decod.pc_q_o\[9\] _02054_ u_decod.pc_q_o\[10\] VGND VGND VPWR VPWR _02149_
+ sky130_fd_sc_hd__a21oi_1
X_05918_ _01207_ VGND VGND VPWR VPWR _01208_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_120_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ u_decod.pc0_q_i\[17\] _01150_ VGND VGND VPWR VPWR _01154_ sky130_fd_sc_hd__or2_1
X_08637_ u_rf.reg29_q\[22\] _03217_ _03291_ u_rf.reg11_q\[22\] VGND VGND VPWR VPWR
+ _03819_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_87_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08568_ u_rf.reg28_q\[19\] _03331_ _03333_ u_rf.reg2_q\[19\] VGND VGND VPWR VPWR
+ _03753_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07519_ u_rf.reg0_q\[22\] _01663_ _01616_ u_rf.reg31_q\[22\] VGND VGND VPWR VPWR
+ _02745_ sky130_fd_sc_hd__a22o_1
X_08499_ _03681_ _03683_ _03685_ _03687_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10530_ _04770_ u_rf.reg15_q\[23\] _05100_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10461_ _05067_ VGND VGND VPWR VPWR _00470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ clknet_leaf_17_clk _00237_ net289 VGND VGND VPWR VPWR u_rf.reg7_q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10392_ _04768_ u_rf.reg13_q\[22\] _05028_ VGND VGND VPWR VPWR _05031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12131_ clknet_leaf_108_clk _00168_ net312 VGND VGND VPWR VPWR u_rf.reg5_q\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12062_ clknet_leaf_1_clk _00099_ net209 VGND VGND VPWR VPWR u_rf.reg3_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_11013_ u_rf.reg22_q\[25\] _04991_ _05355_ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ clknet_leaf_107_clk _01001_ net315 VGND VGND VPWR VPWR u_rf.reg31_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11915_ clknet_leaf_102_clk u_decod.rs1_data\[3\] net336 VGND VGND VPWR VPWR u_decod.rs1_data_q\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_12895_ clknet_leaf_131_clk _00932_ net227 VGND VGND VPWR VPWR u_rf.reg29_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_127 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11846_ clknet_leaf_111_clk _00073_ net317 VGND VGND VPWR VPWR u_rf.reg0_q\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ clknet_leaf_87_clk net160 net362 VGND VGND VPWR VPWR u_decod.pc0_q_i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10728_ _05209_ VGND VGND VPWR VPWR _00595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10659_ u_rf.reg17_q\[19\] _04978_ _05163_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12329_ clknet_leaf_56_clk _00366_ net286 VGND VGND VPWR VPWR u_rf.reg11_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07870_ _03041_ _03042_ _01897_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__o21ai_1
X_06821_ u_rf.reg7_q\[8\] _01559_ _01604_ u_rf.reg3_q\[8\] VGND VGND VPWR VPWR _02075_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06752_ _01059_ _02008_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__nand2_1
X_09540_ _04543_ VGND VGND VPWR VPWR _00073_ sky130_fd_sc_hd__clkbuf_1
X_09471_ _04506_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06683_ u_decod.dec0.funct7\[0\] _01530_ _01549_ u_decod.rf_ff_res_data_i\[5\] _01942_
+ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__a221o_1
X_08422_ u_rf.reg30_q\[12\] _03341_ _03342_ u_rf.reg10_q\[12\] _03613_ VGND VGND VPWR
+ VPWR _03614_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08353_ u_rf.reg30_q\[9\] _03281_ _03283_ u_rf.reg10_q\[9\] _03547_ VGND VGND VPWR
+ VPWR _03548_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07304_ _02446_ _02538_ _01057_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__a21oi_1
X_08284_ u_rf.reg7_q\[6\] _03314_ _03315_ u_rf.reg25_q\[6\] _03481_ VGND VGND VPWR
+ VPWR _03482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07235_ u_rf.reg0_q\[16\] _01662_ _01635_ u_rf.reg9_q\[16\] _02472_ VGND VGND VPWR
+ VPWR _02473_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07166_ _02289_ _02406_ _01688_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06117_ u_decod.rs1_data_q\[16\] VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__buf_4
X_07097_ _02142_ _02339_ _01457_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06048_ _01314_ _01316_ _01317_ _01318_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout222 net223 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_2
XFILLER_0_10_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout211 net220 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout244 net246 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout233 net254 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_2
Xfanout255 net374 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_4
Xfanout299 net301 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_2
Xfanout277 net279 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_4
X_07999_ _03181_ u_decod.dec0.instr_i\[18\] VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__nor2_2
Xfanout266 net270 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_4
Xfanout288 net290 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_4
X_09807_ _04688_ VGND VGND VPWR VPWR _00195_ sky130_fd_sc_hd__clkbuf_1
X_09738_ _04651_ VGND VGND VPWR VPWR _00163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09669_ _04613_ VGND VGND VPWR VPWR _00132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11700_ u_decod.branch_imm_q_o\[28\] _03020_ _05717_ VGND VGND VPWR VPWR _05725_
+ sky130_fd_sc_hd__mux2_1
X_12680_ clknet_leaf_19_clk _00717_ net282 VGND VGND VPWR VPWR u_rf.reg22_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11631_ _04780_ u_rf.reg31_q\[28\] _05679_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11562_ _05651_ VGND VGND VPWR VPWR _00987_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10513_ _04753_ u_rf.reg15_q\[15\] _05089_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11493_ _04778_ u_rf.reg29_q\[27\] _05607_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10444_ _05058_ VGND VGND VPWR VPWR _00462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10375_ _04751_ u_rf.reg13_q\[14\] _05017_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__mux2_1
X_12114_ clknet_leaf_46_clk _00151_ net298 VGND VGND VPWR VPWR u_rf.reg4_q\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ clknet_leaf_64_clk u_decod.exe_ff_res_data_i\[25\] net346 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[25\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_148_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_54_clk _00984_ net303 VGND VGND VPWR VPWR u_rf.reg30_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_160 u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12878_ clknet_leaf_9_clk _00915_ net226 VGND VGND VPWR VPWR u_rf.reg28_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_171 u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 _03320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_182 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11829_ clknet_leaf_115_clk net17 net323 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07020_ _02259_ _02261_ _02263_ _02265_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__or4_1
XFILLER_0_12_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08971_ _04101_ _04123_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__nor2_1
X_07922_ _01268_ _02244_ _01820_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__o21a_1
X_07853_ u_rf.reg24_q\[29\] _01784_ _01668_ u_rf.reg8_q\[29\] VGND VGND VPWR VPWR
+ _03065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06804_ _01332_ _01336_ _01340_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__o21ai_1
X_07784_ u_decod.pc_q_o\[27\] u_decod.pc_q_o\[28\] _02909_ VGND VGND VPWR VPWR _02999_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_97_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ u_rf.reg0_q\[1\] _04430_ _04533_ VGND VGND VPWR VPWR _04535_ sky130_fd_sc_hd__mux2_1
X_06735_ _01328_ _01947_ _01329_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_148_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06666_ u_rf.reg28_q\[5\] _01624_ _01665_ u_rf.reg8_q\[5\] VGND VGND VPWR VPWR _01926_
+ sky130_fd_sc_hd__a22o_1
X_09454_ u_rf.reg1_q\[1\] _04430_ _04496_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08405_ u_rf.reg1_q\[11\] _03446_ _03447_ u_rf.reg14_q\[11\] VGND VGND VPWR VPWR
+ _03598_ sky130_fd_sc_hd__a22o_1
X_09385_ u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__buf_2
X_08336_ u_rf.reg28_q\[8\] _03330_ _03332_ u_rf.reg2_q\[8\] VGND VGND VPWR VPWR _03532_
+ sky130_fd_sc_hd__a22o_1
X_06597_ _01321_ _01324_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08267_ _03459_ _03461_ _03463_ _03465_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_140_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_140_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08198_ u_rf.reg4_q\[2\] _03224_ _03225_ u_rf.reg17_q\[2\] VGND VGND VPWR VPWR _03400_
+ sky130_fd_sc_hd__a22o_1
X_07218_ _01688_ _02350_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07149_ u_decod.dec0.funct3\[2\] _01208_ _02256_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_131_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10160_ _04891_ VGND VGND VPWR VPWR _00345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10091_ u_rf.reg9_q\[25\] _04480_ _04849_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10993_ _05350_ VGND VGND VPWR VPWR _00719_ sky130_fd_sc_hd__clkbuf_1
X_12801_ clknet_leaf_95_clk _00838_ net325 VGND VGND VPWR VPWR u_rf.reg26_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12732_ clknet_leaf_127_clk _00769_ net237 VGND VGND VPWR VPWR u_rf.reg24_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12663_ clknet_leaf_71_clk _00700_ net353 VGND VGND VPWR VPWR u_rf.reg21_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12594_ clknet_leaf_38_clk _00631_ net274 VGND VGND VPWR VPWR u_rf.reg19_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11614_ _05656_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_13_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11545_ _05642_ VGND VGND VPWR VPWR _00979_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_131_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_131_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11476_ _04761_ u_rf.reg29_q\[19\] _05596_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10427_ _05049_ VGND VGND VPWR VPWR _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10358_ _04734_ u_rf.reg13_q\[6\] _05006_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10289_ u_decod.rf_ff_res_data_i\[14\] VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12028_ clknet_leaf_112_clk u_decod.exe_ff_res_data_i\[8\] net321 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_665 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06520_ u_rf.reg25_q\[2\] _01783_ _01784_ u_rf.reg24_q\[2\] _01785_ VGND VGND VPWR
+ VPWR _01786_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_66_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06451_ u_rf.reg6_q\[1\] _01555_ _01580_ u_rf.reg30_q\[1\] _01718_ VGND VGND VPWR
+ VPWR _01719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09170_ u_decod.pc_q_o\[16\] u_decod.branch_imm_q_o\[16\] VGND VGND VPWR VPWR _04296_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06382_ _01651_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_32_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08121_ _03324_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_122_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_122_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08052_ _03178_ _03255_ _03257_ net436 VGND VGND VPWR VPWR u_decod.rs1_data\[31\]
+ sky130_fd_sc_hd__a22o_1
X_07003_ _02249_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_610 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08954_ _01376_ u_decod.branch_imm_q_o\[19\] u_decod.branch_imm_q_o\[18\] _01384_
+ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_110_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07905_ u_rf.reg5_q\[30\] _02664_ _01610_ u_rf.reg12_q\[30\] VGND VGND VPWR VPWR
+ _03115_ sky130_fd_sc_hd__a22o_1
X_08885_ _04048_ _04049_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__nor2_1
X_07836_ _03010_ _03048_ _02723_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_16_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07767_ u_rf.reg16_q\[27\] _02307_ _02379_ u_rf.reg17_q\[27\] VGND VGND VPWR VPWR
+ _02983_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09506_ u_rf.reg1_q\[26\] _04482_ _04518_ VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06718_ u_rf.reg16_q\[6\] _01564_ _01673_ u_rf.reg2_q\[6\] _01975_ VGND VGND VPWR
+ VPWR _01976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07698_ u_decod.rs1_data_q\[26\] _01384_ _01302_ u_decod.rs1_data_q\[2\] _01469_
+ _01466_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__mux4_1
X_09437_ u_decod.rf_ff_res_data_i\[28\] VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_406 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06649_ _01686_ _01909_ _01450_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09368_ _04439_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09299_ _04396_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08319_ u_rf.reg16_q\[7\] _03450_ _03515_ u_rf.reg5_q\[7\] VGND VGND VPWR VPWR _03516_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_113_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_113_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_93 _05463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11330_ _04751_ u_rf.reg27_q\[14\] _05524_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux2_1
XANTENNA_82 _04874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_71 _04544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_60 _03373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ _05492_ VGND VGND VPWR VPWR _00845_ sky130_fd_sc_hd__clkbuf_1
X_13000_ clknet_leaf_92_clk _01037_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[13\]
+ sky130_fd_sc_hd__dfxtp_2
X_11192_ u_rf.reg25_q\[13\] _04966_ _05452_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__mux2_1
X_10212_ _04919_ VGND VGND VPWR VPWR _00369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10143_ _04882_ VGND VGND VPWR VPWR _00337_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10074_ u_rf.reg9_q\[17\] _04463_ _04838_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10976_ _05341_ VGND VGND VPWR VPWR _00711_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12715_ clknet_leaf_136_clk _00752_ net207 VGND VGND VPWR VPWR u_rf.reg23_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12646_ clknet_leaf_3_clk _00683_ net211 VGND VGND VPWR VPWR u_rf.reg21_q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_104_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12577_ clknet_leaf_117_clk _00614_ net326 VGND VGND VPWR VPWR u_rf.reg19_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11528_ _04745_ u_rf.reg30_q\[11\] _05632_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11459_ _05597_ VGND VGND VPWR VPWR _00938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05951_ u_decod.dec0.instr_i\[5\] _01086_ VGND VGND VPWR VPWR _01231_ sky130_fd_sc_hd__nand2_1
X_08670_ u_rf.reg0_q\[23\] _03175_ _03328_ u_rf.reg12_q\[23\] VGND VGND VPWR VPWR
+ _03851_ sky130_fd_sc_hd__a22o_1
X_05882_ _01177_ _01144_ _01178_ VGND VGND VPWR VPWR _01179_ sky130_fd_sc_hd__and3b_1
XFILLER_0_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07621_ u_rf.reg24_q\[24\] _01784_ _02379_ u_rf.reg17_q\[24\] _02842_ VGND VGND VPWR
+ VPWR _02843_ sky130_fd_sc_hd__a221o_1
X_07552_ _02618_ _02776_ _02621_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_37_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06503_ _01313_ _01769_ VGND VGND VPWR VPWR _01770_ sky130_fd_sc_hd__and2b_1
X_07483_ u_rf.reg26_q\[21\] _01642_ _01644_ u_rf.reg20_q\[21\] VGND VGND VPWR VPWR
+ _02711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09222_ u_decod.pc_q_o\[24\] u_decod.branch_imm_q_o\[24\] VGND VGND VPWR VPWR _04340_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06434_ _01494_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__buf_2
XFILLER_0_146_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09153_ _04071_ _04274_ _04275_ _04281_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[13\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06365_ _01634_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08104_ u_rf.reg6_q\[0\] _03305_ _03307_ u_rf.reg13_q\[0\] VGND VGND VPWR VPWR _03308_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09084_ u_decod.pc_q_o\[4\] u_decod.branch_imm_q_o\[4\] VGND VGND VPWR VPWR _04222_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_79_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06296_ _01520_ u_decod.dec0.instr_i\[21\] VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__nor2_2
XFILLER_0_32_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput80 reset_adr_i[23] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_1
XFILLER_0_102_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput91 reset_adr_i[4] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
X_08035_ _03171_ _03172_ _03198_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__and3_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09986_ u_rf.reg8_q\[8\] _04444_ _04790_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux2_1
X_08937_ _01384_ u_decod.branch_imm_q_o\[18\] VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08868_ u_decod.rs1_data_q\[8\] u_decod.branch_imm_q_o\[8\] VGND VGND VPWR VPWR _04035_
+ sky130_fd_sc_hd__nor2_1
X_07819_ u_rf.reg3_q\[28\] _02363_ _01668_ u_rf.reg8_q\[28\] _03032_ VGND VGND VPWR
+ VPWR _03033_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_4_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08799_ _03964_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_123_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10830_ u_rf.reg20_q\[3\] _04945_ _05260_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__mux2_1
X_10761_ _05227_ VGND VGND VPWR VPWR _00610_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_348 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_523 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12500_ clknet_leaf_32_clk _00537_ net263 VGND VGND VPWR VPWR u_rf.reg16_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10692_ u_rf.reg18_q\[2\] _04943_ _05188_ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12431_ clknet_leaf_37_clk _00468_ net273 VGND VGND VPWR VPWR u_rf.reg14_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12362_ clknet_leaf_29_clk _00399_ net257 VGND VGND VPWR VPWR u_rf.reg12_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11313_ _04734_ u_rf.reg27_q\[6\] _05513_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__mux2_1
X_12293_ clknet_leaf_120_clk _00330_ net248 VGND VGND VPWR VPWR u_rf.reg10_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11244_ _05483_ VGND VGND VPWR VPWR _00837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ u_rf.reg25_q\[5\] _04949_ _05441_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10126_ _04873_ VGND VGND VPWR VPWR _00329_ sky130_fd_sc_hd__clkbuf_1
X_10057_ u_rf.reg9_q\[9\] _04446_ _04827_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10959_ _04682_ _04645_ _05295_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__and3_4
XFILLER_0_85_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12629_ clknet_leaf_45_clk _00666_ net298 VGND VGND VPWR VPWR u_rf.reg20_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_06150_ _01394_ _01408_ _01418_ _01419_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__nand4_2
XFILLER_0_79_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06081_ _01291_ _01290_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__nor2_1
Xhold116 u_decod.pc0_q_i\[0\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold105 u_decod.dec0.instr_i\[10\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 u_exe.pc_data_q\[17\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 u_rf.reg19_q\[14\] VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 u_decod.rf_ff_res_data_i\[4\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_74_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09840_ _04705_ VGND VGND VPWR VPWR _00211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09771_ _04668_ VGND VGND VPWR VPWR _00179_ sky130_fd_sc_hd__clkbuf_1
X_06983_ _02225_ _02230_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[11\] sky130_fd_sc_hd__xnor2_1
X_08722_ u_rf.reg26_q\[26\] _03343_ _03285_ u_rf.reg21_q\[26\] VGND VGND VPWR VPWR
+ _03900_ sky130_fd_sc_hd__a22o_1
X_05934_ _01218_ VGND VGND VPWR VPWR u_decod.dec0.rd_o\[4\] sky130_fd_sc_hd__clkbuf_1
X_05865_ u_decod.pc0_q_i\[21\] _01162_ VGND VGND VPWR VPWR _01166_ sky130_fd_sc_hd__nand2_1
X_08653_ u_decod.exe_ff_res_data_i\[22\] _03381_ _03834_ VGND VGND VPWR VPWR _03835_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_1_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05796_ u_decod.pc0_q_i\[2\] u_decod.pc0_q_i\[3\] u_decod.pc0_q_i\[4\] u_decod.pc0_q_i\[5\]
+ VGND VGND VPWR VPWR _01113_ sky130_fd_sc_hd__and4_1
XFILLER_0_89_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08584_ u_rf.reg15_q\[19\] _03301_ _03303_ u_rf.reg24_q\[19\] _03768_ VGND VGND VPWR
+ VPWR _03769_ sky130_fd_sc_hd__a221o_1
X_07604_ _01267_ _01498_ _02136_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07535_ u_rf.reg18_q\[22\] _01787_ _02652_ u_rf.reg23_q\[22\] _02760_ VGND VGND VPWR
+ VPWR _02761_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07466_ _02675_ _02676_ _02694_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09205_ _04318_ _04320_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06417_ _01388_ _01683_ u_decod.rs1_data_q\[8\] u_decod.rs1_data_q\[24\] _01446_
+ _01685_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07397_ _01820_ _02627_ _01365_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_72_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ _04264_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06348_ u_rf.reg3_q\[0\] _01606_ _01610_ u_rf.reg12_q\[0\] _01617_ VGND VGND VPWR
+ VPWR _01618_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_20_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09067_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06279_ _01548_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08018_ _03170_ _03172_ _03205_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__and3_4
XFILLER_0_102_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09969_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12980_ clknet_leaf_23_clk _01017_ net285 VGND VGND VPWR VPWR u_rf.reg31_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11931_ clknet_leaf_86_clk u_decod.rs1_data\[19\] net338 VGND VGND VPWR VPWR u_decod.rs1_data_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_11862_ clknet_leaf_33_clk _00089_ net269 VGND VGND VPWR VPWR u_rf.reg0_q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10813_ _05254_ VGND VGND VPWR VPWR _00635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11793_ clknet_leaf_79_clk net146 net371 VGND VGND VPWR VPWR u_decod.pc0_q_i\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10744_ u_rf.reg18_q\[27\] _04995_ _05210_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10675_ _05181_ VGND VGND VPWR VPWR _00570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12414_ clknet_leaf_123_clk _00451_ net243 VGND VGND VPWR VPWR u_rf.reg14_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12345_ clknet_leaf_57_clk _00382_ net293 VGND VGND VPWR VPWR u_rf.reg11_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_37 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12276_ clknet_leaf_34_clk _00313_ net267 VGND VGND VPWR VPWR u_rf.reg9_q\[25\] sky130_fd_sc_hd__dfrtp_1
X_11227_ u_rf.reg25_q\[30\] _05001_ _05440_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11158_ _05437_ VGND VGND VPWR VPWR _00797_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10109_ u_rf.reg10_q\[1\] _04430_ _04863_ VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__mux2_1
X_11089_ _04782_ u_rf.reg23_q\[29\] _05391_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07320_ u_rf.reg0_q\[18\] _01662_ _01635_ u_rf.reg9_q\[18\] VGND VGND VPWR VPWR _02554_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07251_ _01897_ _02488_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07182_ u_rf.reg7_q\[15\] _01561_ _01642_ u_rf.reg26_q\[15\] VGND VGND VPWR VPWR
+ _02422_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06202_ _01470_ _01471_ _01472_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_367 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06133_ u_decod.rs2_data_q\[19\] _01376_ _01385_ _01402_ _01403_ VGND VGND VPWR VPWR
+ _01404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_395 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06064_ u_decod.rs2_data_q\[7\] u_decod.rs1_data_q\[7\] VGND VGND VPWR VPWR _01335_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_6_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09823_ u_rf.reg6_q\[11\] _04451_ _04695_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ u_rf.reg18_q\[11\] _01591_ _01649_ u_rf.reg4_q\[11\] VGND VGND VPWR VPWR
+ _02214_ sky130_fd_sc_hd__a22o_1
X_09754_ u_rf.reg5_q\[11\] _04451_ _04658_ VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__mux2_1
X_08705_ _03877_ _03879_ _03881_ _03883_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or4_1
X_06897_ net34 _02047_ _02049_ net51 _02051_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__a221o_1
X_09685_ u_rf.reg4_q\[12\] _04453_ _04619_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__mux2_1
X_05917_ _01205_ _01206_ VGND VGND VPWR VPWR _01207_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08636_ u_rf.reg16_q\[22\] _03323_ _03295_ u_rf.reg20_q\[22\] _03817_ VGND VGND VPWR
+ VPWR _03818_ sky130_fd_sc_hd__a221o_1
X_05848_ u_decod.pc0_q_i\[17\] _01150_ VGND VGND VPWR VPWR _01153_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_87_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_139_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05779_ _01100_ VGND VGND VPWR VPWR _01101_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_763 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08567_ net469 _03565_ _03752_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[18\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ u_rf.reg27_q\[15\] _03319_ _03321_ u_rf.reg19_q\[15\] _03686_ VGND VGND VPWR
+ VPWR _03687_ sky130_fd_sc_hd__a221o_1
X_07518_ u_decod.dec0.instr_i\[22\] _01206_ _02646_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07449_ u_decod.pc_q_o\[21\] _02638_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10460_ _04768_ u_rf.reg14_q\[22\] _05064_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ _04250_ _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10391_ _05030_ VGND VGND VPWR VPWR _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12130_ clknet_leaf_131_clk _00167_ net229 VGND VGND VPWR VPWR u_rf.reg5_q\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_131_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12061_ clknet_leaf_119_clk _00098_ net250 VGND VGND VPWR VPWR u_rf.reg3_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11012_ _05360_ VGND VGND VPWR VPWR _00728_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12963_ clknet_leaf_107_clk _01000_ net315 VGND VGND VPWR VPWR u_rf.reg31_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_84_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11914_ clknet_leaf_97_clk u_decod.rs1_data\[2\] net332 VGND VGND VPWR VPWR u_decod.rs1_data_q\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12894_ clknet_leaf_12_clk _00931_ net221 VGND VGND VPWR VPWR u_rf.reg29_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11845_ clknet_leaf_108_clk _00072_ net314 VGND VGND VPWR VPWR u_rf.reg0_q\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ clknet_leaf_89_clk net159 net361 VGND VGND VPWR VPWR u_decod.pc0_q_i\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_126_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10727_ u_rf.reg18_q\[19\] _04978_ _05199_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10658_ _05172_ VGND VGND VPWR VPWR _00562_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10589_ u_rf.reg16_q\[18\] _04976_ _05127_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12328_ clknet_leaf_56_clk _00365_ net291 VGND VGND VPWR VPWR u_rf.reg11_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_584 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12259_ clknet_leaf_108_clk _00296_ net312 VGND VGND VPWR VPWR u_rf.reg9_q\[8\] sky130_fd_sc_hd__dfrtp_1
X_06820_ u_rf.reg5_q\[8\] _01567_ _01593_ u_rf.reg19_q\[8\] _02073_ VGND VGND VPWR
+ VPWR _02074_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06751_ net62 _01487_ _01488_ net48 _02007_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_75_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
X_06682_ _01932_ _01941_ _01678_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__o21a_1
X_09470_ u_rf.reg1_q\[9\] _04446_ _04496_ VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08421_ u_rf.reg26_q\[12\] _03284_ _03345_ u_rf.reg21_q\[12\] VGND VGND VPWR VPWR
+ _03613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_903 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08352_ u_rf.reg26_q\[9\] _03343_ _03286_ u_rf.reg21_q\[9\] VGND VGND VPWR VPWR _03547_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07303_ net100 net42 VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__nand2_1
X_08283_ u_rf.reg1_q\[6\] _03310_ _03312_ u_rf.reg14_q\[6\] VGND VGND VPWR VPWR _03481_
+ sky130_fd_sc_hd__a22o_1
X_07234_ u_rf.reg19_q\[16\] _01594_ _01649_ u_rf.reg4_q\[16\] VGND VGND VPWR VPWR
+ _02472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07165_ _02192_ _02405_ _01451_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06116_ _01385_ _01386_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__nand2_1
X_07096_ _01955_ _02338_ _01685_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06047_ u_decod.rs1_data_q\[1\] _01315_ VGND VGND VPWR VPWR _01318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout212 net220 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_2
Xfanout223 net255 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout256 net257 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_4
Xfanout245 net246 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_4
Xfanout234 net238 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout278 net279 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_4
Xfanout267 net269 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07998_ u_decod.dec0.instr_i\[15\] _03190_ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__and2_2
Xfanout289 net290 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09806_ u_rf.reg6_q\[3\] _04434_ _04684_ VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__mux2_1
X_09737_ u_rf.reg5_q\[3\] _04434_ _04647_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__mux2_1
X_06949_ _01904_ _02001_ _02094_ _02197_ _01475_ _01905_ VGND VGND VPWR VPWR _02198_
+ sky130_fd_sc_hd__mux4_2
Xclkbuf_leaf_66_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09668_ u_rf.reg4_q\[4\] _04436_ _04608_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08619_ u_rf.reg30_q\[21\] _03341_ _03342_ u_rf.reg10_q\[21\] _03801_ VGND VGND VPWR
+ VPWR _03802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09599_ u_rf.reg3_q\[4\] _04436_ _04571_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__mux2_1
X_11630_ _05687_ VGND VGND VPWR VPWR _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11561_ _04778_ u_rf.reg30_q\[27\] _05643_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10512_ _05094_ VGND VGND VPWR VPWR _00494_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_276 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11492_ _05614_ VGND VGND VPWR VPWR _00954_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10443_ _04751_ u_rf.reg14_q\[14\] _05053_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10374_ _05021_ VGND VGND VPWR VPWR _00429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12113_ clknet_leaf_55_clk _00150_ net296 VGND VGND VPWR VPWR u_rf.reg4_q\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_53_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12044_ clknet_leaf_74_clk u_decod.exe_ff_res_data_i\[24\] net356 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[24\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_148_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_57_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_153_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12946_ clknet_leaf_46_clk _00983_ net299 VGND VGND VPWR VPWR u_rf.reg30_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12877_ clknet_leaf_10_clk _00914_ net224 VGND VGND VPWR VPWR u_rf.reg28_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_161 u_decod.dec0.funct7\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_150 _03337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _04911_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 u_decod.rs1_data_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11828_ clknet_leaf_115_clk net16 net328 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_183 net334 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11759_ clknet_leaf_28_clk _00051_ net256 VGND VGND VPWR VPWR u_rf.reg1_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_747 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08970_ _04119_ _04122_ VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__xnor2_1
X_07921_ _01268_ _01269_ _03128_ _03129_ _02332_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__o311a_1
X_07852_ u_rf.reg5_q\[29\] _02664_ _02368_ u_rf.reg26_q\[29\] _03063_ VGND VGND VPWR
+ VPWR _03064_ sky130_fd_sc_hd__a221o_1
Xinput1 icache_instr_i[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_06803_ _01058_ _02052_ _02057_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_leaf_48_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
X_07783_ u_decod.pc_q_o\[27\] _02909_ u_decod.pc_q_o\[28\] VGND VGND VPWR VPWR _02998_
+ sky130_fd_sc_hd__a21oi_1
X_09522_ _04534_ VGND VGND VPWR VPWR _00064_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06734_ _01990_ _01991_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[6\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09453_ _04497_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__clkbuf_1
X_06665_ u_rf.reg24_q\[5\] _01621_ _01649_ u_rf.reg4_q\[5\] _01924_ VGND VGND VPWR
+ VPWR _01925_ sky130_fd_sc_hd__a221o_1
X_09384_ _04450_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08404_ u_rf.reg15_q\[11\] _03373_ _03374_ u_rf.reg24_q\[11\] _03596_ VGND VGND VPWR
+ VPWR _03597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08335_ _03524_ _03526_ _03528_ _03530_ VGND VGND VPWR VPWR _03531_ sky130_fd_sc_hd__or4_1
X_06596_ _01323_ _01763_ _01857_ _01858_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_74_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08266_ u_rf.reg11_q\[5\] _03291_ _03263_ u_rf.reg23_q\[5\] _03464_ VGND VGND VPWR
+ VPWR _03465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08197_ u_rf.reg8_q\[2\] _03216_ _03272_ u_rf.reg29_q\[2\] _03398_ VGND VGND VPWR
+ VPWR _03399_ sky130_fd_sc_hd__a221o_1
X_07217_ _02238_ _02455_ _01464_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07148_ _02374_ _02389_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_89_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07079_ u_rf.reg29_q\[13\] _01627_ _01652_ u_rf.reg22_q\[13\] VGND VGND VPWR VPWR
+ _02323_ sky130_fd_sc_hd__a22o_1
X_10090_ _04854_ VGND VGND VPWR VPWR _00312_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_39_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_98_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12800_ clknet_leaf_114_clk _00837_ net330 VGND VGND VPWR VPWR u_rf.reg26_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ u_rf.reg22_q\[15\] _04970_ _05344_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12731_ clknet_leaf_11_clk _00768_ net222 VGND VGND VPWR VPWR u_rf.reg24_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_12662_ clknet_leaf_49_clk _00699_ net308 VGND VGND VPWR VPWR u_rf.reg21_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_908 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11613_ _05678_ VGND VGND VPWR VPWR _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12593_ clknet_leaf_56_clk _00630_ net286 VGND VGND VPWR VPWR u_rf.reg19_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_703 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11544_ _04761_ u_rf.reg30_q\[19\] _05632_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11475_ _05605_ VGND VGND VPWR VPWR _00946_ sky130_fd_sc_hd__clkbuf_1
X_10426_ _04734_ u_rf.reg14_q\[6\] _05042_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10357_ _05012_ VGND VGND VPWR VPWR _00421_ sky130_fd_sc_hd__clkbuf_1
X_10288_ _04967_ VGND VGND VPWR VPWR _00397_ sky130_fd_sc_hd__clkbuf_1
X_12027_ clknet_leaf_113_clk u_decod.exe_ff_res_data_i\[7\] net322 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12929_ clknet_leaf_95_clk _00966_ net327 VGND VGND VPWR VPWR u_rf.reg30_q\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06450_ u_rf.reg16_q\[1\] _01564_ _01652_ u_rf.reg22_q\[1\] VGND VGND VPWR VPWR _01718_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_574 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06381_ _01572_ _01551_ _01553_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__and3_4
XFILLER_0_126_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08120_ _03249_ VGND VGND VPWR VPWR _03324_ sky130_fd_sc_hd__buf_8
XFILLER_0_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08051_ _03256_ VGND VGND VPWR VPWR _03257_ sky130_fd_sc_hd__buf_2
XFILLER_0_113_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_622 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07002_ _02043_ _02248_ _01457_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _04106_ _04107_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07904_ _03107_ _03109_ _03111_ _03113_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08884_ _01302_ u_decod.branch_imm_q_o\[10\] VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07835_ _01477_ _02960_ _01502_ VGND VGND VPWR VPWR _03048_ sky130_fd_sc_hd__a21boi_1
X_07766_ _02975_ _02977_ _02979_ _02981_ VGND VGND VPWR VPWR _02982_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09505_ _04524_ VGND VGND VPWR VPWR _00057_ sky130_fd_sc_hd__clkbuf_1
X_06717_ u_rf.reg23_q\[6\] _01611_ _01638_ u_rf.reg21_q\[6\] VGND VGND VPWR VPWR _01975_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09436_ _04485_ VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07697_ _02332_ _02911_ _02913_ _02915_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06648_ _01363_ _01683_ _01297_ u_decod.rs1_data_q\[28\] _01446_ _01685_ VGND VGND
+ VPWR VPWR _01909_ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09367_ u_rf.reg2_q\[5\] _04438_ _04428_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__mux2_1
X_06579_ u_rf.reg11_q\[3\] _01583_ _01659_ u_rf.reg14_q\[3\] _01842_ VGND VGND VPWR
+ VPWR _01843_ sky130_fd_sc_hd__a221o_1
X_08318_ _03324_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__buf_8
XANTENNA_50 _03325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09298_ _04385_ u_decod.rs2_data_q\[12\] _04386_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_83 _04981_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _03378_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_72 _04544_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08249_ u_rf.reg7_q\[4\] _03428_ _03429_ u_rf.reg25_q\[4\] _03448_ VGND VGND VPWR
+ VPWR _03449_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 _05463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11260_ u_rf.reg26_q\[13\] u_decod.rf_ff_res_data_i\[13\] _05488_ VGND VGND VPWR
+ VPWR _05492_ sky130_fd_sc_hd__mux2_1
X_10211_ _04757_ u_rf.reg11_q\[17\] _04911_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__mux2_1
X_11191_ _05455_ VGND VGND VPWR VPWR _00812_ sky130_fd_sc_hd__clkbuf_1
X_10142_ u_rf.reg10_q\[17\] _04463_ _04874_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__mux2_1
Xoutput190 net190 VGND VGND VPWR VPWR store_data_o[30] sky130_fd_sc_hd__buf_4
X_10073_ _04845_ VGND VGND VPWR VPWR _00304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_145_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12714_ clknet_leaf_30_clk _00751_ net262 VGND VGND VPWR VPWR u_rf.reg23_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_839 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10975_ u_rf.reg22_q\[7\] _04953_ _05333_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ clknet_leaf_116_clk _00682_ net324 VGND VGND VPWR VPWR u_rf.reg21_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12576_ clknet_leaf_116_clk _00613_ net324 VGND VGND VPWR VPWR u_rf.reg19_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11527_ _05633_ VGND VGND VPWR VPWR _00970_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11458_ _04742_ u_rf.reg29_q\[10\] _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__mux2_1
X_10409_ _05039_ VGND VGND VPWR VPWR _00446_ sky130_fd_sc_hd__clkbuf_1
X_11389_ _05548_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05950_ _01230_ VGND VGND VPWR VPWR u_decod.dec0.unit_o\[3\] sky130_fd_sc_hd__clkbuf_1
X_05881_ u_decod.pc0_q_i\[23\] u_decod.pc0_q_i\[24\] _01168_ u_decod.pc0_q_i\[25\]
+ VGND VGND VPWR VPWR _01178_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07620_ u_rf.reg26_q\[24\] _02368_ _02385_ u_rf.reg20_q\[24\] VGND VGND VPWR VPWR
+ _02842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07551_ _02619_ net48 VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06502_ _01317_ _01435_ _01436_ _01319_ _01432_ VGND VGND VPWR VPWR _01769_ sky130_fd_sc_hd__a221o_1
X_07482_ u_rf.reg0_q\[21\] _01663_ _01601_ u_rf.reg15_q\[21\] _02709_ VGND VGND VPWR
+ VPWR _02710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09221_ _04128_ _04274_ _04275_ _04339_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[23\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_118_215 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06433_ _01445_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09152_ _04278_ _04280_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_831 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06364_ _01513_ _01566_ _01573_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__and3_2
X_08103_ _03306_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__buf_8
XFILLER_0_17_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06295_ _01564_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_8
X_09083_ u_decod.pc_q_o\[4\] u_decod.branch_imm_q_o\[4\] VGND VGND VPWR VPWR _04221_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_79_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput81 reset_adr_i[24] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_1
XFILLER_0_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput70 reset_adr_i[14] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
X_08034_ u_rf.reg6_q\[31\] _03235_ _03236_ u_rf.reg13_q\[31\] _03239_ VGND VGND VPWR
+ VPWR _03240_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput92 reset_adr_i[5] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_92_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09985_ _04798_ VGND VGND VPWR VPWR _00263_ sky130_fd_sc_hd__clkbuf_1
X_08936_ _04042_ _04093_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__nor2_1
X_08867_ _03998_ _04034_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__nor2_1
X_07818_ u_rf.reg5_q\[28\] _02664_ _02360_ u_rf.reg9_q\[28\] VGND VGND VPWR VPWR _03032_
+ sky130_fd_sc_hd__a22o_1
X_08798_ _03966_ _03968_ _03970_ _03972_ VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_123_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07749_ _02919_ _02965_ _01481_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10760_ u_rf.reg19_q\[2\] _04943_ _05224_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09419_ u_decod.rf_ff_res_data_i\[22\] VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10691_ _05190_ VGND VGND VPWR VPWR _00577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12430_ clknet_leaf_27_clk _00467_ net258 VGND VGND VPWR VPWR u_rf.reg14_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12361_ clknet_leaf_21_clk _00398_ net280 VGND VGND VPWR VPWR u_rf.reg12_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11312_ _05519_ VGND VGND VPWR VPWR _00869_ sky130_fd_sc_hd__clkbuf_1
X_12292_ clknet_leaf_107_clk _00329_ net314 VGND VGND VPWR VPWR u_rf.reg10_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_11243_ u_rf.reg26_q\[5\] u_decod.rf_ff_res_data_i\[5\] _05477_ VGND VGND VPWR VPWR
+ _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11174_ _05446_ VGND VGND VPWR VPWR _00804_ sky130_fd_sc_hd__clkbuf_1
X_10125_ u_rf.reg10_q\[9\] _04446_ _04863_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__mux2_1
X_10056_ _04836_ VGND VGND VPWR VPWR _00296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10958_ _05331_ VGND VGND VPWR VPWR _00703_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12628_ clknet_leaf_34_clk _00665_ net268 VGND VGND VPWR VPWR u_rf.reg20_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10889_ _05294_ VGND VGND VPWR VPWR _00671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12559_ clknet_leaf_35_clk _00596_ net275 VGND VGND VPWR VPWR u_rf.reg18_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold106 u_exe.pc_data_q\[2\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06080_ _01300_ _01304_ _01346_ _01347_ _01350_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__o311a_2
Xhold117 u_decod.rf_ff_res_data_i\[3\] VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_111_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold139 u_exe.pc_data_q\[3\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 u_decod.dec0.instr_i\[11\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ u_rf.reg5_q\[19\] _04467_ _04658_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__mux2_1
X_06982_ _02089_ _02227_ _02229_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__a21o_1
X_08721_ u_rf.reg8_q\[26\] _03407_ _03408_ u_rf.reg29_q\[26\] _03898_ VGND VGND VPWR
+ VPWR _03899_ sky130_fd_sc_hd__a221o_1
X_05933_ net502 u_decod.dec0.rd_v VGND VGND VPWR VPWR _01218_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08652_ u_decod.rf_ff_res_data_i\[22\] _03382_ _03833_ _03404_ VGND VGND VPWR VPWR
+ _03834_ sky130_fd_sc_hd__a22o_1
X_05864_ u_decod.pc0_q_i\[21\] _01162_ VGND VGND VPWR VPWR _01165_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_750 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07603_ _01425_ _02787_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_1_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05795_ net516 _01105_ _01101_ net91 _01112_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__a221o_4
X_08583_ u_rf.reg6_q\[19\] _03387_ _03388_ u_rf.reg13_q\[19\] VGND VGND VPWR VPWR
+ _03768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07534_ u_rf.reg24_q\[22\] _01622_ _01780_ u_rf.reg29_q\[22\] VGND VGND VPWR VPWR
+ _02760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07465_ _01485_ _02677_ _02678_ _02693_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09204_ _04323_ _04324_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__or2b_1
XFILLER_0_107_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06416_ _01684_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07396_ _01763_ _02244_ _01395_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09135_ _04265_ _04260_ _04257_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__o21a_1
XFILLER_0_60_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06347_ u_rf.reg23_q\[0\] _01613_ _01616_ u_rf.reg31_q\[0\] VGND VGND VPWR VPWR _01617_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09066_ u_decod.instr_operation_q\[5\] _01485_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__nand2_4
XFILLER_0_72_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06278_ _01517_ _01527_ _01547_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_20_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08017_ _03188_ _03209_ _03205_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__and3_4
XFILLER_0_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09968_ _04423_ _04788_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_125_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08919_ _01289_ u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__nor2_1
X_11930_ clknet_leaf_101_clk u_decod.rs1_data\[18\] net338 VGND VGND VPWR VPWR u_decod.rs1_data_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_09899_ u_decod.rf_ff_res_data_i\[10\] VGND VGND VPWR VPWR _04742_ sky130_fd_sc_hd__buf_2
X_11861_ clknet_leaf_66_clk _00088_ net355 VGND VGND VPWR VPWR u_rf.reg0_q\[24\] sky130_fd_sc_hd__dfrtp_1
X_10812_ u_rf.reg19_q\[27\] _04995_ _05246_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__mux2_1
X_11792_ clknet_leaf_79_clk net144 net371 VGND VGND VPWR VPWR u_decod.pc0_q_i\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10743_ _05217_ VGND VGND VPWR VPWR _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10674_ u_rf.reg17_q\[26\] _04993_ _05174_ VGND VGND VPWR VPWR _05181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12413_ clknet_leaf_13_clk _00450_ net245 VGND VGND VPWR VPWR u_rf.reg14_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12344_ clknet_leaf_63_clk _00381_ net342 VGND VGND VPWR VPWR u_rf.reg11_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12275_ clknet_leaf_54_clk _00312_ net302 VGND VGND VPWR VPWR u_rf.reg9_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11226_ _05473_ VGND VGND VPWR VPWR _00829_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_56_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ u_rf.reg24_q\[29\] _04999_ _05427_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10108_ _04864_ VGND VGND VPWR VPWR _00320_ sky130_fd_sc_hd__clkbuf_1
X_11088_ _05400_ VGND VGND VPWR VPWR _00764_ sky130_fd_sc_hd__clkbuf_1
X_10039_ u_rf.reg9_q\[0\] _04421_ _04827_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07250_ _02089_ _02487_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07181_ u_rf.reg15_q\[15\] _02371_ _01610_ u_rf.reg12_q\[15\] _02420_ VGND VGND VPWR
+ VPWR _02421_ sky130_fd_sc_hd__a221o_1
X_06201_ _01451_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_379 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06132_ u_decod.rs2_data_q\[18\] _01384_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06063_ _01328_ _01333_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__nor2_1
X_09822_ _04696_ VGND VGND VPWR VPWR _00202_ sky130_fd_sc_hd__clkbuf_1
X_09753_ _04659_ VGND VGND VPWR VPWR _00170_ sky130_fd_sc_hd__clkbuf_1
X_08704_ u_rf.reg31_q\[25\] _03290_ _03292_ u_rf.reg11_q\[25\] _03882_ VGND VGND VPWR
+ VPWR _03883_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _02206_ _02208_ _02210_ _02212_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__or4_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05916_ _01069_ _01080_ _01072_ u_decod.dec0.instr_i\[4\] VGND VGND VPWR VPWR _01206_
+ sky130_fd_sc_hd__and4bb_4
X_09684_ _04621_ VGND VGND VPWR VPWR _00139_ sky130_fd_sc_hd__clkbuf_1
X_06896_ _01478_ _02095_ _02146_ _01505_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__o211a_1
X_08635_ u_rf.reg4_q\[22\] _03264_ _03266_ u_rf.reg17_q\[22\] VGND VGND VPWR VPWR
+ _03817_ sky130_fd_sc_hd__a22o_1
X_05847_ net514 _01142_ _01132_ net72 _01152_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__a221o_2
XTAP_TAPCELL_ROW_87_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ u_decod.exe_ff_res_data_i\[18\] _03381_ _03751_ VGND VGND VPWR VPWR _03752_
+ sky130_fd_sc_hd__a21o_1
X_05778_ u_ifetch.reset_n_q net369 VGND VGND VPWR VPWR _01100_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_138_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07517_ _01773_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08497_ u_rf.reg16_q\[15\] _03323_ _03325_ u_rf.reg5_q\[15\] VGND VGND VPWR VPWR
+ _03686_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_274 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_639 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07448_ u_decod.pc_q_o\[21\] _02638_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07379_ u_rf.reg3_q\[19\] _01605_ _01638_ u_rf.reg21_q\[19\] VGND VGND VPWR VPWR
+ _02611_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09118_ u_decod.pc_q_o\[9\] u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _04251_
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_70_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ _04766_ u_rf.reg13_q\[21\] _05028_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09049_ u_decod.instr_operation_q\[0\] _04188_ u_decod.instr_operation_q\[5\] u_decod.instr_operation_q\[4\]
+ VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12060_ clknet_leaf_128_clk _00097_ net236 VGND VGND VPWR VPWR u_rf.reg3_q\[1\] sky130_fd_sc_hd__dfrtp_1
X_11011_ u_rf.reg22_q\[24\] _04989_ _05355_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ clknet_leaf_129_clk _00999_ net235 VGND VGND VPWR VPWR u_rf.reg31_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12893_ clknet_leaf_16_clk _00930_ net250 VGND VGND VPWR VPWR u_rf.reg29_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_11913_ clknet_leaf_102_clk u_decod.rs1_data\[1\] net336 VGND VGND VPWR VPWR u_decod.rs1_data_q\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_157_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11844_ clknet_leaf_130_clk _00071_ net234 VGND VGND VPWR VPWR u_rf.reg0_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11775_ clknet_leaf_87_clk net156 net360 VGND VGND VPWR VPWR u_decod.pc0_q_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_155_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10726_ _05208_ VGND VGND VPWR VPWR _00594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10657_ u_rf.reg17_q\[18\] _04976_ _05163_ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_508 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10588_ _05135_ VGND VGND VPWR VPWR _00529_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12327_ clknet_leaf_5_clk _00364_ net213 VGND VGND VPWR VPWR u_rf.reg11_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12258_ clknet_leaf_129_clk _00295_ net234 VGND VGND VPWR VPWR u_rf.reg9_q\[7\] sky130_fd_sc_hd__dfrtp_1
X_11209_ u_rf.reg25_q\[21\] _04983_ _05463_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_118_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12189_ clknet_leaf_13_clk _00226_ net245 VGND VGND VPWR VPWR u_rf.reg7_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_06750_ net39 _01489_ _01490_ net57 VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06681_ _01934_ _01936_ _01938_ _01940_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_69_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08420_ u_rf.reg31_q\[12\] _03504_ _03505_ u_rf.reg11_q\[12\] _03611_ VGND VGND VPWR
+ VPWR _03612_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08351_ u_rf.reg8_q\[9\] _03271_ _03273_ u_rf.reg29_q\[9\] _03545_ VGND VGND VPWR
+ VPWR _03546_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08282_ u_rf.reg0_q\[6\] _03176_ _03329_ u_rf.reg12_q\[6\] _03479_ VGND VGND VPWR
+ VPWR _03480_ sky130_fd_sc_hd__a221o_1
X_07302_ _02495_ _02536_ _01425_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07233_ u_rf.reg31_q\[16\] _01615_ _01658_ u_rf.reg14_q\[16\] _02470_ VGND VGND VPWR
+ VPWR _02471_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07164_ _02403_ _02404_ _01460_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06115_ u_decod.rs2_data_q\[18\] _01384_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__nand2_1
X_07095_ u_decod.rs1_data_q\[14\] _01446_ _01753_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06046_ u_decod.rs1_data_q\[2\] u_decod.rs2_data_q\[2\] VGND VGND VPWR VPWR _01317_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_136_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout213 net220 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout202 net204 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_4
Xfanout224 net226 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net253 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_4
Xfanout235 net238 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_4
Xfanout279 net311 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__buf_2
Xfanout268 net269 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_89_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07997_ u_decod.dec0.instr_i\[19\] _03201_ _03199_ VGND VGND VPWR VPWR _03203_ sky130_fd_sc_hd__and3_4
Xfanout257 net260 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_4
X_09805_ _04687_ VGND VGND VPWR VPWR _00194_ sky130_fd_sc_hd__clkbuf_1
X_09736_ _04650_ VGND VGND VPWR VPWR _00162_ sky130_fd_sc_hd__clkbuf_1
X_06948_ _01460_ _01823_ _02196_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__a21o_1
X_09667_ _04612_ VGND VGND VPWR VPWR _00131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08618_ u_rf.reg26_q\[21\] _03284_ _03286_ u_rf.reg21_q\[21\] VGND VGND VPWR VPWR
+ _03801_ sky130_fd_sc_hd__a22o_1
X_06879_ u_decod.dec0.funct7\[4\] _01529_ _01548_ u_decod.rf_ff_res_data_i\[9\] _02130_
+ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09598_ _04575_ VGND VGND VPWR VPWR _00099_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08549_ u_rf.reg7_q\[18\] _03314_ _03388_ u_rf.reg13_q\[18\] _03734_ VGND VGND VPWR
+ VPWR _03735_ sky130_fd_sc_hd__a221o_1
X_11560_ _05650_ VGND VGND VPWR VPWR _00986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10511_ _04751_ u_rf.reg15_q\[14\] _05089_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11491_ _04776_ u_rf.reg29_q\[26\] _05607_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_150_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10442_ _05057_ VGND VGND VPWR VPWR _00461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10373_ _04749_ u_rf.reg13_q\[13\] _05017_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12112_ clknet_leaf_23_clk _00149_ net284 VGND VGND VPWR VPWR u_rf.reg4_q\[21\] sky130_fd_sc_hd__dfrtp_1
X_12043_ clknet_leaf_73_clk u_decod.exe_ff_res_data_i\[23\] net358 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[23\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_53_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ clknet_leaf_54_clk _00982_ net296 VGND VGND VPWR VPWR u_rf.reg30_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_140 _02604_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ clknet_leaf_19_clk _00913_ net281 VGND VGND VPWR VPWR u_rf.reg28_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_151 _03356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 u_decod.rs1_data_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11827_ clknet_leaf_115_clk net15 net328 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_162 u_decod.dec0.funct7\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_195 _04911_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11758_ clknet_leaf_6_clk _00050_ net215 VGND VGND VPWR VPWR u_rf.reg1_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ u_rf.reg18_q\[10\] _04959_ _05199_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11689_ _05719_ VGND VGND VPWR VPWR _01046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_817 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_759 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07920_ _01273_ _03083_ _01270_ _01272_ VGND VGND VPWR VPWR _03129_ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07851_ u_rf.reg0_q\[29\] _01664_ _02385_ u_rf.reg20_q\[29\] VGND VGND VPWR VPWR
+ _03063_ sky130_fd_sc_hd__a22o_1
X_07782_ _02994_ _02997_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[27\] sky130_fd_sc_hd__xnor2_1
Xinput2 icache_instr_i[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_06802_ _01764_ _02053_ _02054_ _02056_ _01339_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__o32a_1
XFILLER_0_79_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09521_ u_rf.reg0_q\[0\] _04421_ _04533_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__mux2_1
X_06733_ _01744_ _01944_ _01946_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_84_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ u_rf.reg1_q\[0\] _04421_ _04496_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__mux2_1
X_06664_ u_rf.reg30_q\[5\] _01578_ _01599_ u_rf.reg15_q\[5\] VGND VGND VPWR VPWR _01924_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09383_ u_rf.reg2_q\[10\] _04448_ _04449_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__mux2_1
X_08403_ u_rf.reg6_q\[11\] _03305_ _03307_ u_rf.reg13_q\[11\] VGND VGND VPWR VPWR
+ _03596_ sky130_fd_sc_hd__a22o_1
X_06595_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] u_decod.pc_q_o\[4\] _01764_ VGND
+ VGND VPWR VPWR _01858_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08334_ u_rf.reg31_q\[8\] _03290_ _03292_ u_rf.reg11_q\[8\] _03529_ VGND VGND VPWR
+ VPWR _03530_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08265_ u_rf.reg22_q\[5\] _03274_ _03276_ u_rf.reg3_q\[5\] VGND VGND VPWR VPWR _03464_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_115_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08196_ u_rf.reg22_q\[2\] _03218_ _03219_ u_rf.reg3_q\[2\] VGND VGND VPWR VPWR _03398_
+ sky130_fd_sc_hd__a22o_1
X_07216_ _01267_ _01467_ _02136_ _02454_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_144_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07147_ _02378_ _02382_ _02384_ _02388_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07078_ u_rf.reg11_q\[13\] _01584_ _01598_ u_rf.reg13_q\[13\] _02321_ VGND VGND VPWR
+ VPWR _02322_ sky130_fd_sc_hd__a221o_1
X_06029_ u_decod.rs2_data_q\[11\] u_decod.rs1_data_q\[11\] VGND VGND VPWR VPWR _01300_
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_153_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09719_ _04639_ VGND VGND VPWR VPWR _00156_ sky130_fd_sc_hd__clkbuf_1
X_10991_ _05349_ VGND VGND VPWR VPWR _00718_ sky130_fd_sc_hd__clkbuf_1
X_12730_ clknet_leaf_64_clk _00767_ net341 VGND VGND VPWR VPWR u_rf.reg23_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12661_ clknet_leaf_47_clk _00698_ net301 VGND VGND VPWR VPWR u_rf.reg21_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11612_ _04761_ u_rf.reg31_q\[19\] _05668_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12592_ clknet_leaf_31_clk _00629_ net263 VGND VGND VPWR VPWR u_rf.reg19_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11543_ _05641_ VGND VGND VPWR VPWR _00978_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11474_ _04759_ u_rf.reg29_q\[18\] _05596_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10425_ _05048_ VGND VGND VPWR VPWR _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10356_ _04732_ u_rf.reg13_q\[5\] _05006_ VGND VGND VPWR VPWR _05012_ sky130_fd_sc_hd__mux2_1
X_10287_ u_rf.reg12_q\[13\] _04966_ _04960_ VGND VGND VPWR VPWR _04967_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12026_ clknet_leaf_97_clk u_decod.exe_ff_res_data_i\[6\] net331 VGND VGND VPWR VPWR
+ u_decod.rf_ff_res_data_i\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12928_ clknet_leaf_115_clk _00965_ net323 VGND VGND VPWR VPWR u_rf.reg30_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12859_ clknet_leaf_13_clk _00896_ net242 VGND VGND VPWR VPWR u_rf.reg28_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06380_ _01649_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__buf_6
XFILLER_0_126_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_311 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08050_ u_decod.dec0.instr_i\[5\] _01224_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07001_ _01864_ _02247_ _01684_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08952_ _01363_ u_decod.branch_imm_q_o\[20\] VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_110_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07903_ u_rf.reg31_q\[30\] _01777_ _02380_ u_rf.reg10_q\[30\] _03112_ VGND VGND VPWR
+ VPWR _03113_ sky130_fd_sc_hd__a221o_1
X_08883_ _01302_ u_decod.branch_imm_q_o\[10\] VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__nor2_1
X_07834_ u_decod.instr_operation_q\[3\] _01263_ _01432_ _01414_ _03046_ VGND VGND
+ VPWR VPWR _03047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07765_ u_rf.reg9_q\[27\] _02360_ _01668_ u_rf.reg8_q\[27\] _02980_ VGND VGND VPWR
+ VPWR _02981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09504_ u_rf.reg1_q\[25\] _04480_ _04518_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__mux2_1
X_07696_ _02781_ _01409_ _02914_ _01284_ VGND VGND VPWR VPWR _02915_ sky130_fd_sc_hd__a22o_1
X_06716_ u_rf.reg7_q\[6\] _01560_ _01641_ u_rf.reg26_q\[6\] _01973_ VGND VGND VPWR
+ VPWR _01974_ sky130_fd_sc_hd__a221o_1
X_09435_ u_rf.reg2_q\[27\] _04484_ _04470_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06647_ _01505_ _01907_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_577 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09366_ u_decod.rf_ff_res_data_i\[5\] VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__buf_2
X_06578_ u_rf.reg19_q\[3\] _01594_ _01652_ u_rf.reg22_q\[3\] VGND VGND VPWR VPWR _01842_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_40 _03285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09297_ _04395_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08317_ u_rf.reg7_q\[7\] _03428_ _03429_ u_rf.reg25_q\[7\] _03513_ VGND VGND VPWR
+ VPWR _03514_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_62 _03388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _03331_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _05006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08248_ u_rf.reg1_q\[4\] _03446_ _03447_ u_rf.reg14_q\[4\] VGND VGND VPWR VPWR _03448_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_73 _04647_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 _05512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08179_ _03187_ VGND VGND VPWR VPWR _03381_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10210_ _04918_ VGND VGND VPWR VPWR _00368_ sky130_fd_sc_hd__clkbuf_1
X_11190_ u_rf.reg25_q\[12\] _04964_ _05452_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__mux2_1
X_10141_ _04881_ VGND VGND VPWR VPWR _00336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput191 net191 VGND VGND VPWR VPWR store_data_o[31] sky130_fd_sc_hd__buf_4
Xoutput180 net180 VGND VGND VPWR VPWR store_data_o[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10072_ u_rf.reg9_q\[16\] _04461_ _04838_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10974_ _05340_ VGND VGND VPWR VPWR _00710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12713_ clknet_leaf_22_clk _00750_ net284 VGND VGND VPWR VPWR u_rf.reg23_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12644_ clknet_leaf_112_clk _00681_ net321 VGND VGND VPWR VPWR u_rf.reg21_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12575_ clknet_leaf_137_clk _00612_ net205 VGND VGND VPWR VPWR u_rf.reg19_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11526_ _04742_ u_rf.reg30_q\[10\] _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11457_ _05584_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__buf_8
XFILLER_0_68_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10408_ _04784_ u_rf.reg13_q\[30\] _05005_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11388_ _05559_ VGND VGND VPWR VPWR _00905_ sky130_fd_sc_hd__clkbuf_1
X_10339_ u_rf.reg12_q\[30\] _05001_ _04938_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__mux2_1
X_12009_ clknet_leaf_80_clk u_exe.bu_pc_res\[22\] net371 VGND VGND VPWR VPWR u_exe.pc_data_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_05880_ u_decod.pc0_q_i\[24\] u_decod.pc0_q_i\[25\] _01171_ VGND VGND VPWR VPWR _01177_
+ sky130_fd_sc_hd__and3_4
X_07550_ _02773_ _01485_ _02774_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__and3b_1
XFILLER_0_108_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06501_ _01317_ _01763_ _01764_ u_decod.pc_q_o\[2\] _01767_ VGND VGND VPWR VPWR _01768_
+ sky130_fd_sc_hd__o221ai_1
X_09220_ _04337_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__xnor2_1
X_07481_ u_rf.reg7_q\[21\] _01561_ _01605_ u_rf.reg3_q\[21\] VGND VGND VPWR VPWR _02709_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_227 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06432_ _01694_ _01436_ _01695_ _01700_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09151_ _04279_ _04272_ _04269_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06363_ u_rf.reg24_q\[0\] _01622_ _01625_ u_rf.reg28_q\[0\] _01632_ VGND VGND VPWR
+ VPWR _01633_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08102_ _03236_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__buf_8
X_09082_ _04197_ _04218_ _04219_ _04220_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[3\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08033_ u_rf.reg15_q\[31\] _03237_ _03238_ u_rf.reg24_q\[31\] VGND VGND VPWR VPWR
+ _03239_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06294_ _01563_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__buf_6
XFILLER_0_32_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput82 reset_adr_i[25] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_1
Xinput71 reset_adr_i[15] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
XFILLER_0_130_904 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput60 load_data_i[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XFILLER_0_142_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput93 reset_adr_i[6] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09984_ u_rf.reg8_q\[7\] _04442_ _04790_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08935_ _04091_ _04092_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__xor2_1
X_08866_ _04032_ _04033_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__xnor2_1
X_07817_ u_rf.reg23_q\[28\] _02652_ _01654_ u_rf.reg22_q\[28\] _03030_ VGND VGND VPWR
+ VPWR _03031_ sky130_fd_sc_hd__a221o_1
X_08797_ u_rf.reg22_q\[29\] _03275_ _03366_ u_rf.reg19_q\[29\] _03971_ VGND VGND VPWR
+ VPWR _03972_ sky130_fd_sc_hd__a221o_1
X_07748_ _02684_ _02778_ _02874_ _02964_ _01476_ _02685_ VGND VGND VPWR VPWR _02965_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_140_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07679_ u_rf.reg16_q\[25\] _01564_ _01636_ u_rf.reg9_q\[25\] _02898_ VGND VGND VPWR
+ VPWR _02899_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09418_ _04473_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_158 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10690_ u_rf.reg18_q\[1\] _04941_ _05188_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09349_ _01531_ _01536_ _04425_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_43_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12360_ clknet_leaf_59_clk _00397_ net289 VGND VGND VPWR VPWR u_rf.reg12_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11311_ _04732_ u_rf.reg27_q\[5\] _05513_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12291_ clknet_leaf_107_clk _00328_ net314 VGND VGND VPWR VPWR u_rf.reg10_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11242_ _05482_ VGND VGND VPWR VPWR _00836_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11173_ u_rf.reg25_q\[4\] _04947_ _05441_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10124_ _04872_ VGND VGND VPWR VPWR _00328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10055_ u_rf.reg9_q\[8\] _04444_ _04827_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10957_ u_rf.reg21_q\[31\] _05003_ _05296_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_51_clk _00664_ net303 VGND VGND VPWR VPWR u_rf.reg20_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ u_rf.reg20_q\[31\] _05003_ _05259_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12558_ clknet_leaf_28_clk _00595_ net256 VGND VGND VPWR VPWR u_rf.reg18_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 u_exe.pc_data_q\[22\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ clknet_leaf_25_clk _00526_ net270 VGND VGND VPWR VPWR u_rf.reg16_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11509_ _04726_ u_rf.reg30_q\[2\] _05621_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_228 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold118 u_exe.pc_data_q\[0\] VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 u_decod.rf_ff_res_data_i\[0\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_1
XFILLER_0_110_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _01079_ _01250_ _01243_ _02228_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__a211oi_4
X_08720_ u_rf.reg22_q\[26\] _03409_ _03410_ u_rf.reg3_q\[26\] VGND VGND VPWR VPWR
+ _03898_ sky130_fd_sc_hd__a22o_1
X_05932_ _01217_ VGND VGND VPWR VPWR u_decod.dec0.rd_o\[3\] sky130_fd_sc_hd__clkbuf_1
X_05863_ net498 _01142_ _01132_ net77 _01164_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__a221o_1
X_08651_ _03823_ _03832_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__or2_1
X_07602_ _01437_ _02821_ _02822_ _02824_ _01279_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_1_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05794_ _01110_ _01106_ _01111_ VGND VGND VPWR VPWR _01112_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08582_ u_rf.reg1_q\[19\] _03311_ _03313_ u_rf.reg14_q\[19\] _03766_ VGND VGND VPWR
+ VPWR _03767_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07533_ u_rf.reg17_q\[22\] _02379_ _02380_ u_rf.reg10_q\[22\] _02758_ VGND VGND VPWR
+ VPWR _02759_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_637 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07464_ _01443_ _02683_ _02690_ _02692_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09203_ u_decod.pc_q_o\[21\] u_decod.branch_imm_q_o\[21\] VGND VGND VPWR VPWR _04324_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06415_ u_decod.rs2_data_q\[3\] VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__inv_2
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09134_ _04258_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__inv_2
X_07395_ _02581_ _02625_ _01424_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06346_ _01615_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_8
X_09065_ _01063_ _04200_ _04197_ _04205_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[1\]
+ sky130_fd_sc_hd__a22o_1
X_06277_ _01531_ _01522_ _01533_ _01546_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08016_ _03188_ _03173_ _03199_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__and3_4
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09967_ u_decod.rf_ff_rd_adr_q_i\[0\] _04424_ _01531_ _01535_ VGND VGND VPWR VPWR
+ _04788_ sky130_fd_sc_hd__or4_4
X_08918_ _04042_ _04078_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_125_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _04741_ VGND VGND VPWR VPWR _00233_ sky130_fd_sc_hd__clkbuf_1
X_08849_ u_decod.rs1_data_q\[5\] u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _04019_
+ sky130_fd_sc_hd__and2_1
X_11860_ clknet_leaf_38_clk _00087_ net277 VGND VGND VPWR VPWR u_rf.reg0_q\[23\] sky130_fd_sc_hd__dfrtp_1
X_10811_ _05253_ VGND VGND VPWR VPWR _00634_ sky130_fd_sc_hd__clkbuf_1
X_11791_ clknet_leaf_79_clk net143 net371 VGND VGND VPWR VPWR u_decod.pc0_q_i\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10742_ u_rf.reg18_q\[26\] _04993_ _05210_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10673_ _05180_ VGND VGND VPWR VPWR _00569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12412_ clknet_leaf_128_clk _00449_ net236 VGND VGND VPWR VPWR u_rf.reg14_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12343_ clknet_leaf_49_clk _00380_ net352 VGND VGND VPWR VPWR u_rf.reg11_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_153_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12274_ clknet_leaf_41_clk _00311_ net278 VGND VGND VPWR VPWR u_rf.reg9_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11225_ u_rf.reg25_q\[29\] _04999_ _05463_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ _05436_ VGND VGND VPWR VPWR _00796_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11087_ _04780_ u_rf.reg23_q\[28\] _05391_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__mux2_1
X_10107_ u_rf.reg10_q\[0\] _04421_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__mux2_1
X_10038_ _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11989_ clknet_leaf_89_clk u_exe.bu_pc_res\[2\] net361 VGND VGND VPWR VPWR u_exe.pc_data_q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06200_ u_decod.rs1_data_q\[4\] _01297_ _01363_ u_decod.rs1_data_q\[28\] _01460_
+ _01461_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07180_ u_rf.reg25_q\[15\] _01783_ _02419_ u_rf.reg28_q\[15\] VGND VGND VPWR VPWR
+ _02420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06131_ _01381_ _01400_ _01401_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06062_ _01310_ _01323_ _01309_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09821_ u_rf.reg6_q\[10\] _04448_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__mux2_1
X_09752_ u_rf.reg5_q\[10\] _04448_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08703_ u_rf.reg9_q\[25\] _03294_ _03296_ u_rf.reg20_q\[25\] VGND VGND VPWR VPWR
+ _03882_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ u_rf.reg7_q\[11\] _01561_ _01595_ u_rf.reg19_q\[11\] _02211_ VGND VGND VPWR
+ VPWR _02212_ sky130_fd_sc_hd__a221o_1
X_05915_ _01072_ _01070_ VGND VGND VPWR VPWR _01205_ sky130_fd_sc_hd__nor2_1
X_09683_ u_rf.reg4_q\[11\] _04451_ _04619_ VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__mux2_1
X_06895_ _01493_ _02044_ _02145_ u_decod.rs2_data_q\[0\] VGND VGND VPWR VPWR _02146_
+ sky130_fd_sc_hd__a211o_1
X_05846_ _01150_ _01144_ _01151_ VGND VGND VPWR VPWR _01152_ sky130_fd_sc_hd__and3b_1
X_08634_ u_rf.reg9_q\[22\] _03348_ _03300_ u_rf.reg15_q\[22\] _03815_ VGND VGND VPWR
+ VPWR _03816_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_87_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05777_ _01098_ VGND VGND VPWR VPWR _01099_ sky130_fd_sc_hd__buf_4
X_08565_ u_decod.rf_ff_res_data_i\[18\] _03382_ _03750_ _03404_ VGND VGND VPWR VPWR
+ _03751_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07516_ _02742_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[22\] sky130_fd_sc_hd__buf_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08496_ u_rf.reg0_q\[15\] _03420_ _03421_ u_rf.reg12_q\[15\] _03684_ VGND VGND VPWR
+ VPWR _03685_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07447_ _01364_ _01361_ _02637_ _02332_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__o31a_1
XFILLER_0_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07378_ u_rf.reg18_q\[19\] _01592_ _01650_ u_rf.reg4_q\[19\] _02609_ VGND VGND VPWR
+ VPWR _02610_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09117_ u_decod.pc_q_o\[9\] u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _04250_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06329_ _01513_ _01558_ _01577_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__and3_2
XFILLER_0_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09048_ _04177_ _04187_ _02781_ VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_142_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11010_ _05359_ VGND VGND VPWR VPWR _00727_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ clknet_leaf_118_clk _00998_ net326 VGND VGND VPWR VPWR u_rf.reg31_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_51_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ clknet_leaf_99_clk u_decod.rs1_data\[0\] net330 VGND VGND VPWR VPWR u_decod.rs1_data_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12892_ clknet_leaf_128_clk _00929_ net236 VGND VGND VPWR VPWR u_rf.reg29_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11843_ clknet_leaf_119_clk _00070_ net250 VGND VGND VPWR VPWR u_rf.reg0_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11774_ clknet_leaf_87_clk net145 net360 VGND VGND VPWR VPWR u_decod.pc0_q_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_155_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10725_ u_rf.reg18_q\[18\] _04976_ _05199_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__mux2_1
X_10656_ _05171_ VGND VGND VPWR VPWR _00561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10587_ u_rf.reg16_q\[17\] _04974_ _05127_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12326_ clknet_leaf_138_clk _00363_ net210 VGND VGND VPWR VPWR u_rf.reg11_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12257_ clknet_leaf_17_clk _00294_ net251 VGND VGND VPWR VPWR u_rf.reg9_q\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11208_ _05464_ VGND VGND VPWR VPWR _00820_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12188_ clknet_leaf_127_clk _00225_ net237 VGND VGND VPWR VPWR u_rf.reg7_q\[1\] sky130_fd_sc_hd__dfrtp_1
X_11139_ u_rf.reg24_q\[20\] _04980_ _05427_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06680_ u_rf.reg10_q\[5\] _01656_ _01652_ u_rf.reg22_q\[5\] _01939_ VGND VGND VPWR
+ VPWR _01940_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08350_ u_rf.reg22_q\[9\] _03275_ _03277_ u_rf.reg3_q\[9\] VGND VGND VPWR VPWR _03545_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07301_ _02456_ _02535_ _01757_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08281_ u_rf.reg28_q\[6\] _03331_ _03333_ u_rf.reg2_q\[6\] VGND VGND VPWR VPWR _03479_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07232_ u_rf.reg7_q\[16\] _01560_ _01641_ u_rf.reg26_q\[16\] VGND VGND VPWR VPWR
+ _02470_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_640 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07163_ u_decod.rs1_data_q\[30\] _01454_ _02136_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06114_ u_decod.rs2_data_q\[18\] _01384_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07094_ _02334_ _02335_ _02336_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06045_ u_decod.rs1_data_q\[1\] _01315_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_130_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout214 net220 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_2
Xfanout203 net204 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_4
Xfanout225 net226 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
X_09804_ u_rf.reg6_q\[2\] _04432_ _04684_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__mux2_1
Xfanout247 net248 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout236 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_4
Xfanout269 net270 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07996_ _03171_ _03201_ _03199_ VGND VGND VPWR VPWR _03202_ sky130_fd_sc_hd__and3_4
Xfanout258 net260 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09735_ u_rf.reg5_q\[2\] _04432_ _04647_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__mux2_1
X_06947_ u_decod.rs1_data_q\[11\] _01454_ _01685_ _02136_ VGND VGND VPWR VPWR _02196_
+ sky130_fd_sc_hd__o211a_1
X_09666_ u_rf.reg4_q\[3\] _04434_ _04608_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__mux2_1
X_08617_ u_rf.reg31_q\[21\] _03504_ _03505_ u_rf.reg11_q\[21\] _03799_ VGND VGND VPWR
+ VPWR _03800_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06878_ _02120_ _02129_ _01678_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05829_ _01099_ _01136_ _01137_ _01138_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__a31o_1
XFILLER_0_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09597_ u_rf.reg3_q\[3\] _04434_ _04571_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__mux2_1
X_08548_ u_rf.reg30_q\[18\] _03200_ _03285_ u_rf.reg21_q\[18\] VGND VGND VPWR VPWR
+ _03734_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_137_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ u_decod.pc0_q_i\[14\] _03565_ _03668_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[14\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11490_ _05613_ VGND VGND VPWR VPWR _00953_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10510_ _05093_ VGND VGND VPWR VPWR _00493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10441_ _04749_ u_rf.reg14_q\[13\] _05053_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_150_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10372_ _05020_ VGND VGND VPWR VPWR _00428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12111_ clknet_leaf_42_clk _00148_ net275 VGND VGND VPWR VPWR u_rf.reg4_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12042_ clknet_leaf_65_clk u_decod.exe_ff_res_data_i\[22\] net346 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[22\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_53_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_148_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ clknet_leaf_55_clk _00981_ net285 VGND VGND VPWR VPWR u_rf.reg30_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_152 _03366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 _03202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 _01615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12875_ clknet_leaf_2_clk _00912_ net223 VGND VGND VPWR VPWR u_rf.reg28_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_163 u_decod.exe_ff_res_data_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11826_ clknet_leaf_115_clk net14 net328 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_174 u_rf.reg2_q\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 net441 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11757_ clknet_leaf_25_clk _00049_ net280 VGND VGND VPWR VPWR u_rf.reg1_q\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_196 _05017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_134_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_134_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10708_ _05187_ VGND VGND VPWR VPWR _05199_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_64_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11688_ u_decod.branch_imm_q_o\[22\] _02744_ _05717_ VGND VGND VPWR VPWR _05719_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10639_ _05162_ VGND VGND VPWR VPWR _00553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12309_ clknet_leaf_54_clk _00346_ net296 VGND VGND VPWR VPWR u_rf.reg10_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07850_ u_rf.reg13_q\[29\] _02376_ _01777_ u_rf.reg31_q\[29\] _03061_ VGND VGND VPWR
+ VPWR _03062_ sky130_fd_sc_hd__a221o_1
X_07781_ _02229_ _02996_ VGND VGND VPWR VPWR _02997_ sky130_fd_sc_hd__nor2_1
X_06801_ _01307_ _01763_ _01819_ _02055_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__o211a_1
X_09520_ _04532_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__buf_8
X_06732_ _01713_ u_decod.exe_ff_res_data_i\[6\] _01989_ VGND VGND VPWR VPWR _01990_
+ sky130_fd_sc_hd__a21o_1
Xinput3 icache_instr_i[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09451_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__buf_6
X_06663_ _01923_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[5\] sky130_fd_sc_hd__inv_2
XFILLER_0_87_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09382_ _04427_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__buf_6
XFILLER_0_59_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08402_ _03588_ _03590_ _03592_ _03594_ VGND VGND VPWR VPWR _03595_ sky130_fd_sc_hd__or4_1
X_06594_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] u_decod.pc_q_o\[4\] VGND VGND VPWR
+ VPWR _01857_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08333_ u_rf.reg9_q\[8\] _03294_ _03296_ u_rf.reg20_q\[8\] VGND VGND VPWR VPWR _03529_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_125_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_125_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_145_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08264_ u_rf.reg16_q\[5\] _03323_ _03280_ u_rf.reg30_q\[5\] _03462_ VGND VGND VPWR
+ VPWR _03463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08195_ u_rf.reg31_q\[2\] _03289_ _03291_ u_rf.reg11_q\[2\] _03396_ VGND VGND VPWR
+ VPWR _03397_ sky130_fd_sc_hd__a221o_1
X_07215_ _01367_ _01447_ _01685_ _02136_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07146_ u_rf.reg20_q\[14\] _02385_ _02386_ u_rf.reg27_q\[14\] _02387_ VGND VGND VPWR
+ VPWR _02388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07077_ u_rf.reg30_q\[13\] _01579_ _01591_ u_rf.reg18_q\[13\] VGND VGND VPWR VPWR
+ _02321_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06028_ _01296_ _01298_ VGND VGND VPWR VPWR _01299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_668 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09718_ u_rf.reg4_q\[28\] _04486_ _04630_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__mux2_1
X_07979_ _03180_ u_decod.exe_ff_rd_adr_q_i\[0\] u_decod.exe_ff_rd_adr_q_i\[2\] _03181_
+ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o221a_1
X_10990_ u_rf.reg22_q\[14\] _04968_ _05344_ VGND VGND VPWR VPWR _05349_ sky130_fd_sc_hd__mux2_1
X_09649_ u_rf.reg3_q\[28\] _04486_ _04593_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12660_ clknet_leaf_30_clk _00697_ net262 VGND VGND VPWR VPWR u_rf.reg21_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11611_ _05677_ VGND VGND VPWR VPWR _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12591_ clknet_leaf_38_clk _00628_ net274 VGND VGND VPWR VPWR u_rf.reg19_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_116_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_116_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_46_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11542_ _04759_ u_rf.reg30_q\[18\] _05632_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ _05604_ VGND VGND VPWR VPWR _00945_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10424_ _04732_ u_rf.reg14_q\[5\] _05042_ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10355_ _05011_ VGND VGND VPWR VPWR _00420_ sky130_fd_sc_hd__clkbuf_1
X_10286_ u_decod.rf_ff_res_data_i\[13\] VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__buf_2
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12025_ clknet_leaf_98_clk u_decod.exe_ff_res_data_i\[5\] net330 VGND VGND VPWR VPWR
+ u_decod.rf_ff_res_data_i\[5\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12927_ clknet_leaf_131_clk _00964_ net233 VGND VGND VPWR VPWR u_rf.reg30_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12858_ clknet_leaf_61_clk _00895_ net341 VGND VGND VPWR VPWR u_rf.reg27_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11809_ clknet_leaf_106_clk net27 net319 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12789_ clknet_leaf_47_clk _00826_ net301 VGND VGND VPWR VPWR u_rf.reg25_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_107_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_107_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_125_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07000_ u_decod.rs1_data_q\[12\] _01445_ _01494_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08951_ _01363_ u_decod.branch_imm_q_o\[20\] VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_110_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07902_ u_rf.reg7_q\[30\] _01562_ _02363_ u_rf.reg3_q\[30\] VGND VGND VPWR VPWR _03112_
+ sky130_fd_sc_hd__a22o_1
X_08882_ _04042_ _04047_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__nor2_1
X_07833_ u_decod.rs2_data_q\[29\] u_decod.rs1_data_q\[29\] _02781_ VGND VGND VPWR
+ VPWR _03046_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07764_ u_rf.reg30_q\[27\] _01581_ _02419_ u_rf.reg28_q\[27\] VGND VGND VPWR VPWR
+ _02980_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09503_ _04523_ VGND VGND VPWR VPWR _00056_ sky130_fd_sc_hd__clkbuf_1
X_07695_ _01285_ _01435_ _01432_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06715_ u_rf.reg18_q\[6\] _01591_ _01669_ u_rf.reg27_q\[6\] VGND VGND VPWR VPWR _01973_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09434_ u_decod.rf_ff_res_data_i\[27\] VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__buf_2
XFILLER_0_94_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06646_ _01750_ _01825_ _01866_ _01906_ _01478_ _01475_ VGND VGND VPWR VPWR _01907_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09365_ _04437_ VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__clkbuf_1
X_06577_ _01834_ _01836_ _01838_ _01840_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__or4_1
XANTENNA_41 _03290_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_30 _03224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _04385_ u_decod.rs2_data_q\[11\] _04386_ VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_10_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08316_ u_rf.reg1_q\[7\] _03446_ _03447_ u_rf.reg14_q\[7\] VGND VGND VPWR VPWR _03513_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08247_ _03312_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__buf_8
XANTENNA_74 _04764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _03407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_52 _03332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_96 _05535_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _05017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08178_ net441 _03259_ _03380_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[1\]
+ sky130_fd_sc_hd__a22o_1
X_07129_ _01601_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__buf_6
Xoutput170 net170 VGND VGND VPWR VPWR store_data_o[12] sky130_fd_sc_hd__clkbuf_4
X_10140_ u_rf.reg10_q\[16\] _04461_ _04874_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__mux2_1
Xoutput181 net181 VGND VGND VPWR VPWR store_data_o[22] sky130_fd_sc_hd__buf_4
X_10071_ _04844_ VGND VGND VPWR VPWR _00303_ sky130_fd_sc_hd__clkbuf_1
Xoutput192 net192 VGND VGND VPWR VPWR store_data_o[3] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_145_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973_ u_rf.reg22_q\[6\] _04951_ _05333_ VGND VGND VPWR VPWR _05340_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12712_ clknet_leaf_58_clk _00749_ net291 VGND VGND VPWR VPWR u_rf.reg23_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_115 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12643_ clknet_leaf_107_clk _00680_ net315 VGND VGND VPWR VPWR u_rf.reg21_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12574_ clknet_leaf_1_clk _00611_ net221 VGND VGND VPWR VPWR u_rf.reg19_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11525_ _05620_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__buf_8
XFILLER_0_80_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11456_ _05595_ VGND VGND VPWR VPWR _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10407_ _05038_ VGND VGND VPWR VPWR _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11387_ u_rf.reg28_q\[9\] net471 _05549_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__mux2_1
X_10338_ u_decod.rf_ff_res_data_i\[30\] VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__buf_2
X_12008_ clknet_leaf_80_clk u_exe.bu_pc_res\[21\] net371 VGND VGND VPWR VPWR u_exe.pc_data_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10269_ _04954_ VGND VGND VPWR VPWR _00391_ sky130_fd_sc_hd__clkbuf_1
X_07480_ u_rf.reg5_q\[21\] _01569_ _01595_ u_rf.reg19_q\[21\] _02707_ VGND VGND VPWR
+ VPWR _02708_ sky130_fd_sc_hd__a221o_1
X_06500_ _01318_ _01694_ _01765_ _01766_ VGND VGND VPWR VPWR _01767_ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_126 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06431_ _01696_ _01698_ _01699_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__or3_1
X_09150_ _04270_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06362_ u_rf.reg29_q\[0\] _01628_ _01631_ u_rf.reg17_q\[0\] VGND VGND VPWR VPWR _01632_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_716 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08101_ _03304_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__buf_6
X_09081_ _04011_ _04206_ VGND VGND VPWR VPWR _04220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06293_ _01538_ _01514_ _01515_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__and3_2
XFILLER_0_140_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08032_ u_decod.dec0.instr_i\[19\] _03172_ _03201_ VGND VGND VPWR VPWR _03238_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_79_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput72 reset_adr_i[16] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XFILLER_0_130_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput61 load_data_i[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
XFILLER_0_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput50 load_data_i[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
Xinput83 reset_adr_i[26] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
Xinput94 reset_adr_i[7] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09983_ _04797_ VGND VGND VPWR VPWR _00262_ sky130_fd_sc_hd__clkbuf_1
X_08934_ _04086_ _04089_ _04085_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08865_ _04025_ net379 _04024_ VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__a21o_1
X_07816_ u_rf.reg6_q\[28\] _01557_ _02375_ u_rf.reg11_q\[28\] VGND VGND VPWR VPWR
+ _03030_ sky130_fd_sc_hd__a22o_1
X_08796_ u_rf.reg3_q\[29\] _03276_ _03282_ u_rf.reg10_q\[29\] VGND VGND VPWR VPWR
+ _03971_ sky130_fd_sc_hd__a22o_1
X_07747_ u_decod.rs1_data_q\[27\] _01376_ u_decod.rs1_data_q\[11\] u_decod.rs1_data_q\[3\]
+ _01469_ _01466_ VGND VGND VPWR VPWR _02964_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07678_ u_rf.reg0_q\[25\] _01662_ _01666_ u_rf.reg8_q\[25\] VGND VGND VPWR VPWR _02898_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09417_ u_rf.reg2_q\[21\] _04472_ _04470_ VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_619 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06629_ u_rf.reg5_q\[4\] _01569_ _01594_ u_rf.reg19_q\[4\] _01890_ VGND VGND VPWR
+ VPWR _01891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _01534_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11310_ _05518_ VGND VGND VPWR VPWR _00868_ sky130_fd_sc_hd__clkbuf_1
X_09279_ _01427_ VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12290_ clknet_leaf_129_clk _00327_ net234 VGND VGND VPWR VPWR u_rf.reg10_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11241_ u_rf.reg26_q\[4\] net512 _05477_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__mux2_1
X_11172_ _05445_ VGND VGND VPWR VPWR _00803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10123_ u_rf.reg10_q\[8\] _04444_ _04863_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10054_ _04835_ VGND VGND VPWR VPWR _00295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10956_ _05330_ VGND VGND VPWR VPWR _00702_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10887_ _05293_ VGND VGND VPWR VPWR _00670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12626_ clknet_leaf_40_clk _00663_ net278 VGND VGND VPWR VPWR u_rf.reg20_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12557_ clknet_leaf_6_clk _00594_ net216 VGND VGND VPWR VPWR u_rf.reg18_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold108 u_exe.pc_data_q\[5\] VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__dlygate4sd3_1
X_12488_ clknet_leaf_60_clk _00525_ net289 VGND VGND VPWR VPWR u_rf.reg16_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11508_ _05623_ VGND VGND VPWR VPWR _00961_ sky130_fd_sc_hd__clkbuf_1
Xhold119 u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _04724_ u_rf.reg29_q\[1\] _05585_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_74_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _01075_ _01078_ _01084_ _01089_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05931_ net479 u_decod.dec0.rd_v VGND VGND VPWR VPWR _01217_ sky130_fd_sc_hd__and2_1
X_05862_ _01162_ _01144_ _01163_ VGND VGND VPWR VPWR _01164_ sky130_fd_sc_hd__and3b_1
X_08650_ _03825_ _03827_ _03829_ _03831_ VGND VGND VPWR VPWR _03832_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07601_ _01278_ _01435_ _02823_ _01432_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05793_ u_decod.pc0_q_i\[2\] u_decod.pc0_q_i\[3\] u_decod.pc0_q_i\[4\] VGND VGND
+ VPWR VPWR _01111_ sky130_fd_sc_hd__a21o_1
X_08581_ u_rf.reg7_q\[19\] _03369_ _03370_ u_rf.reg25_q\[19\] VGND VGND VPWR VPWR
+ _03766_ sky130_fd_sc_hd__a22o_1
X_07532_ u_rf.reg30_q\[22\] _01580_ _01625_ u_rf.reg28_q\[22\] VGND VGND VPWR VPWR
+ _02758_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_105_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07463_ _02618_ _02691_ _02621_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09202_ u_decod.pc_q_o\[21\] u_decod.branch_imm_q_o\[21\] VGND VGND VPWR VPWR _04323_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_91_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06414_ _01267_ _01430_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__and2_2
X_09133_ _04262_ _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07394_ _02535_ _02624_ _01757_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06345_ _01614_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__buf_6
XFILLER_0_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_231 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09064_ _04198_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__xnor2_1
X_06276_ _01541_ _01543_ _01545_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08015_ u_rf.reg8_q\[31\] _03216_ _03217_ u_rf.reg29_q\[31\] _03220_ VGND VGND VPWR
+ VPWR _03221_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_262 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09966_ _04787_ VGND VGND VPWR VPWR _00255_ sky130_fd_sc_hd__clkbuf_1
X_08917_ _04074_ net383 VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__xnor2_1
X_09897_ _04740_ u_rf.reg7_q\[9\] _04722_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__mux2_1
X_08848_ u_decod.rs1_data_q\[5\] u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _04018_
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_96_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
X_08779_ u_decod.exe_ff_res_data_i\[28\] _03187_ _03382_ u_decod.rf_ff_res_data_i\[28\]
+ _03954_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a221o_1
X_10810_ u_rf.reg19_q\[26\] _04993_ _05246_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__mux2_1
X_11790_ clknet_leaf_83_clk net142 net365 VGND VGND VPWR VPWR u_decod.pc0_q_i\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10741_ _05216_ VGND VGND VPWR VPWR _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10672_ u_rf.reg17_q\[25\] _04991_ _05174_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__mux2_1
X_12411_ clknet_leaf_13_clk _00448_ net243 VGND VGND VPWR VPWR u_rf.reg14_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_20_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_23_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12342_ clknet_leaf_49_clk _00379_ net308 VGND VGND VPWR VPWR u_rf.reg11_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12273_ clknet_leaf_56_clk _00310_ net287 VGND VGND VPWR VPWR u_rf.reg9_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_346 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11224_ _05472_ VGND VGND VPWR VPWR _00828_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ u_rf.reg24_q\[28\] _04997_ _05427_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11086_ _05399_ VGND VGND VPWR VPWR _00763_ sky130_fd_sc_hd__clkbuf_1
X_10106_ _04862_ VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_87_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
X_10037_ _04643_ _04644_ _04825_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__and3_4
XFILLER_0_98_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11988_ clknet_leaf_88_clk u_exe.bu_pc_res\[1\] net360 VGND VGND VPWR VPWR u_exe.pc_data_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ u_rf.reg21_q\[22\] _04985_ _05319_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_693 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12609_ clknet_leaf_118_clk _00646_ net326 VGND VGND VPWR VPWR u_rf.reg20_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_11_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06130_ u_decod.rs2_data_q\[17\] _01380_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__nor2_1
XFILLER_0_152_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06061_ _01311_ _01321_ _01331_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__and3b_1
XFILLER_0_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09820_ _04683_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__buf_6
XFILLER_0_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09751_ _04646_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__buf_8
X_06963_ u_rf.reg16_q\[11\] _01564_ _01583_ u_rf.reg11_q\[11\] VGND VGND VPWR VPWR
+ _02211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_107_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ u_rf.reg30_q\[25\] _03280_ _03282_ u_rf.reg10_q\[25\] _03880_ VGND VGND VPWR
+ VPWR _03881_ sky130_fd_sc_hd__a221o_1
X_05914_ _01092_ _01200_ _01203_ u_decod.dec0.jalr VGND VGND VPWR VPWR _01204_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06894_ _01315_ _02144_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__nor2_1
X_09682_ _04620_ VGND VGND VPWR VPWR _00138_ sky130_fd_sc_hd__clkbuf_1
X_05845_ u_decod.pc0_q_i\[14\] u_decod.pc0_q_i\[15\] net405 u_decod.pc0_q_i\[16\]
+ VGND VGND VPWR VPWR _01151_ sky130_fd_sc_hd__a31o_1
X_08633_ u_rf.reg19_q\[22\] _03247_ _03202_ u_rf.reg10_q\[22\] VGND VGND VPWR VPWR
+ _03815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05776_ u_decod.flush_v net361 VGND VGND VPWR VPWR _01098_ sky130_fd_sc_hd__and2b_1
X_08564_ _03740_ _03749_ VGND VGND VPWR VPWR _03750_ sky130_fd_sc_hd__or2_2
XFILLER_0_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07515_ _02722_ _02730_ _02736_ _02741_ VGND VGND VPWR VPWR _02742_ sky130_fd_sc_hd__or4_1
XFILLER_0_76_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_435 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08495_ u_rf.reg28_q\[15\] _03556_ _03557_ u_rf.reg2_q\[15\] VGND VGND VPWR VPWR
+ _03684_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_60 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07446_ _01395_ _02674_ _01362_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07377_ u_rf.reg6_q\[19\] _01556_ _01653_ u_rf.reg22_q\[19\] VGND VGND VPWR VPWR
+ _02609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06328_ _01597_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_8
X_09116_ _04041_ _04207_ _04208_ _04249_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[8\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09047_ _04176_ _04189_ u_decod.instr_operation_q\[3\] VGND VGND VPWR VPWR _04190_
+ sky130_fd_sc_hd__a21boi_1
X_06259_ _01087_ _01199_ u_decod.dec0.jalr VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__a21o_1
X_09949_ u_decod.rf_ff_res_data_i\[26\] VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_69_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_51_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ clknet_leaf_115_clk _00997_ net324 VGND VGND VPWR VPWR u_rf.reg31_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11911_ clknet_leaf_91_clk u_decod.rs2_data_nxt\[32\] net345 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[32\] sky130_fd_sc_hd__dfrtp_2
X_12891_ clknet_leaf_12_clk _00928_ net221 VGND VGND VPWR VPWR u_rf.reg29_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_11842_ clknet_leaf_119_clk _00069_ net247 VGND VGND VPWR VPWR u_rf.reg0_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11773_ clknet_leaf_87_clk net134 net360 VGND VGND VPWR VPWR u_decod.pc0_q_i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_155_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_827 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10724_ _05207_ VGND VGND VPWR VPWR _00593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10655_ u_rf.reg17_q\[17\] _04974_ _05163_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10586_ _05134_ VGND VGND VPWR VPWR _00528_ sky130_fd_sc_hd__clkbuf_1
X_12325_ clknet_leaf_125_clk _00362_ net240 VGND VGND VPWR VPWR u_rf.reg11_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12256_ clknet_leaf_119_clk _00293_ net248 VGND VGND VPWR VPWR u_rf.reg9_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_11207_ u_rf.reg25_q\[20\] _04980_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12187_ clknet_leaf_13_clk _00224_ net244 VGND VGND VPWR VPWR u_rf.reg7_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_11138_ _05404_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__buf_6
X_11069_ _05390_ VGND VGND VPWR VPWR _00755_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_0_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07300_ _01950_ _02137_ _02346_ _01747_ _01464_ _01468_ VGND VGND VPWR VPWR _02535_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08280_ u_decod.pc0_q_i\[5\] _03259_ _03478_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[5\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07231_ u_rf.reg15_q\[16\] _01600_ _01608_ u_rf.reg12_q\[16\] _02468_ VGND VGND VPWR
+ VPWR _02469_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07162_ _01371_ _01447_ _02136_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06113_ u_decod.rs1_data_q\[18\] VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07093_ u_decod.pc_q_o\[14\] _02284_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_368 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06044_ u_decod.rs2_data_q\[1\] VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_130_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout204 net210 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_130_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout215 net216 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_4
Xfanout226 net255 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout237 net238 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_4
X_09803_ _04686_ VGND VGND VPWR VPWR _00193_ sky130_fd_sc_hd__clkbuf_1
Xfanout259 net260 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_2
X_07995_ u_decod.dec0.instr_i\[17\] _03191_ VGND VGND VPWR VPWR _03201_ sky130_fd_sc_hd__nor2_2
Xfanout248 net252 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_4
X_06946_ _02189_ _02194_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__or2_1
X_09734_ _04649_ VGND VGND VPWR VPWR _00161_ sky130_fd_sc_hd__clkbuf_1
X_09665_ _04611_ VGND VGND VPWR VPWR _00130_ sky130_fd_sc_hd__clkbuf_1
X_06877_ _02122_ _02124_ _02126_ _02128_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__or4_1
X_08616_ u_rf.reg9_q\[21\] _03293_ _03349_ u_rf.reg20_q\[21\] VGND VGND VPWR VPWR
+ _03799_ sky130_fd_sc_hd__a22o_1
X_05828_ net488 _01118_ _01119_ net68 VGND VGND VPWR VPWR _01138_ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09596_ _04574_ VGND VGND VPWR VPWR _00098_ sky130_fd_sc_hd__clkbuf_1
X_08547_ u_rf.reg18_q\[18\] _03352_ _03275_ u_rf.reg22_q\[18\] _03732_ VGND VGND VPWR
+ VPWR _03733_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05759_ u_decod.dec0.funct7\[3\] u_decod.dec0.funct7\[2\] u_decod.dec0.funct7\[4\]
+ _01081_ VGND VGND VPWR VPWR _01082_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_137_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_602 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08478_ u_decod.exe_ff_res_data_i\[14\] _03381_ _03667_ VGND VGND VPWR VPWR _03668_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07429_ u_rf.reg25_q\[20\] _01576_ _01784_ u_rf.reg24_q\[20\] _02658_ VGND VGND VPWR
+ VPWR _02659_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10440_ _05056_ VGND VGND VPWR VPWR _00460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10371_ _04747_ u_rf.reg13_q\[12\] _05017_ VGND VGND VPWR VPWR _05020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ clknet_leaf_28_clk _00147_ net256 VGND VGND VPWR VPWR u_rf.reg4_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12041_ clknet_leaf_65_clk u_decod.exe_ff_res_data_i\[21\] net355 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[21\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_53_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_148_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ clknet_leaf_44_clk _00980_ net295 VGND VGND VPWR VPWR u_rf.reg30_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_120 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12874_ clknet_leaf_26_clk _00911_ net266 VGND VGND VPWR VPWR u_rf.reg28_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_142 _03232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 _01615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_175 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11825_ clknet_leaf_105_clk net13 net321 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_164 u_decod.instr_unit_q\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 _03366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_186 _01468_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11756_ clknet_leaf_12_clk _00048_ net221 VGND VGND VPWR VPWR u_rf.reg1_q\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_197 u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_126_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10707_ _05198_ VGND VGND VPWR VPWR _00585_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11687_ _05718_ VGND VGND VPWR VPWR _01045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_189 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10638_ u_rf.reg17_q\[9\] _04957_ _05152_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_538 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10569_ _05125_ VGND VGND VPWR VPWR _00520_ sky130_fd_sc_hd__clkbuf_1
X_12308_ clknet_leaf_23_clk _00345_ net267 VGND VGND VPWR VPWR u_rf.reg10_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12239_ clknet_leaf_41_clk _00276_ net278 VGND VGND VPWR VPWR u_rf.reg8_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07780_ _02089_ _02487_ _02863_ _02995_ VGND VGND VPWR VPWR _02996_ sky130_fd_sc_hd__and4_1
X_06800_ _01307_ _01434_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__nand2_1
X_06731_ _01679_ _01987_ _01988_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__a21o_1
Xinput4 icache_instr_i[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ _04423_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__nor2_4
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08401_ u_rf.reg30_q\[11\] _03341_ _03342_ u_rf.reg10_q\[11\] _03593_ VGND VGND VPWR
+ VPWR _03594_ sky130_fd_sc_hd__a221o_1
X_06662_ _01901_ _01902_ _01922_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06593_ net59 _01487_ _01488_ net45 _01855_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__a221o_1
X_09381_ u_decod.rf_ff_res_data_i\[10\] VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__buf_2
XFILLER_0_74_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08332_ u_rf.reg30_q\[8\] _03281_ _03283_ u_rf.reg10_q\[8\] _03527_ VGND VGND VPWR
+ VPWR _03528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08263_ u_rf.reg27_q\[5\] _03246_ _03324_ u_rf.reg5_q\[5\] VGND VGND VPWR VPWR _03462_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_49_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07214_ _01820_ _02452_ _01390_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08194_ u_rf.reg9_q\[2\] _03212_ _03213_ u_rf.reg20_q\[2\] VGND VGND VPWR VPWR _03396_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07145_ u_rf.reg23_q\[14\] _01613_ _01622_ u_rf.reg24_q\[14\] VGND VGND VPWR VPWR
+ _02387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07076_ u_rf.reg20_q\[13\] _01645_ _01671_ u_rf.reg27_q\[13\] _02319_ VGND VGND VPWR
+ VPWR _02320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06027_ u_decod.rs2_data_q\[12\] _01297_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_58_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07978_ u_decod.dec0.instr_i\[16\] _01521_ u_decod.exe_ff_rd_adr_q_i\[4\] _03171_
+ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__o22a_1
X_09717_ _04638_ VGND VGND VPWR VPWR _00155_ sky130_fd_sc_hd__clkbuf_1
X_06929_ _01897_ _02178_ _02090_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09648_ _04601_ VGND VGND VPWR VPWR _00123_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09579_ u_rf.reg0_q\[28\] _04486_ _04555_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_67_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12590_ clknet_leaf_7_clk _00627_ net219 VGND VGND VPWR VPWR u_rf.reg19_q\[19\] sky130_fd_sc_hd__dfrtp_1
X_11610_ _04759_ u_rf.reg31_q\[18\] _05668_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11541_ _05640_ VGND VGND VPWR VPWR _00977_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_46_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11472_ _04757_ u_rf.reg29_q\[17\] _05596_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10423_ _05047_ VGND VGND VPWR VPWR _00452_ sky130_fd_sc_hd__clkbuf_1
X_10354_ _04730_ u_rf.reg13_q\[4\] _05006_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_76_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10285_ _04965_ VGND VGND VPWR VPWR _00396_ sky130_fd_sc_hd__clkbuf_1
X_12024_ clknet_leaf_113_clk u_decod.exe_ff_res_data_i\[4\] net322 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12926_ clknet_leaf_133_clk _00963_ net231 VGND VGND VPWR VPWR u_rf.reg30_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_12857_ clknet_leaf_63_clk _00894_ net341 VGND VGND VPWR VPWR u_rf.reg27_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_500 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11808_ clknet_leaf_106_clk net26 net320 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12788_ clknet_leaf_32_clk _00825_ net263 VGND VGND VPWR VPWR u_rf.reg25_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_235 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11739_ clknet_leaf_58_clk _00031_ net343 VGND VGND VPWR VPWR u_rf.reg2_q\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_94_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08950_ _04101_ _04105_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__nor2_1
XFILLER_0_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07901_ u_rf.reg25_q\[30\] _01783_ _01780_ u_rf.reg29_q\[30\] _03110_ VGND VGND VPWR
+ VPWR _03111_ sky130_fd_sc_hd__a221o_1
X_08881_ _04045_ _04046_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__xnor2_1
X_07832_ _01263_ _03044_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07763_ u_rf.reg23_q\[27\] _02652_ _01654_ u_rf.reg22_q\[27\] _02978_ VGND VGND VPWR
+ VPWR _02979_ sky130_fd_sc_hd__a221o_1
X_09502_ u_rf.reg1_q\[24\] _04478_ _04518_ VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07694_ _01277_ _01280_ _02912_ _01411_ _01286_ VGND VGND VPWR VPWR _02913_ sky130_fd_sc_hd__a311o_1
XFILLER_0_78_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06714_ u_rf.reg3_q\[6\] _01605_ _01658_ u_rf.reg14_q\[6\] _01971_ VGND VGND VPWR
+ VPWR _01972_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ _04483_ VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06645_ _01705_ _01904_ _01905_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ u_rf.reg2_q\[4\] _04436_ _04428_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08315_ u_rf.reg15_q\[7\] _03373_ _03374_ u_rf.reg24_q\[7\] _03511_ VGND VGND VPWR
+ VPWR _03512_ sky130_fd_sc_hd__a221o_1
X_06576_ u_rf.reg5_q\[3\] _01569_ _01561_ u_rf.reg7_q\[3\] _01839_ VGND VGND VPWR
+ VPWR _01840_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_20 _01667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_31 _03264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ _04394_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_1
XFILLER_0_145_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08246_ _03310_ VGND VGND VPWR VPWR _03446_ sky130_fd_sc_hd__buf_8
XANTENNA_42 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _04764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_64 _03420_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_53 _03333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 _05100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _05585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08177_ u_decod.exe_ff_res_data_i\[1\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[1\]
+ _03379_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__a221o_1
X_07128_ u_rf.reg31_q\[14\] _01777_ _02367_ u_rf.reg14_q\[14\] _02369_ VGND VGND VPWR
+ VPWR _02370_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_844 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07059_ _02284_ _02285_ _02303_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__o21bai_1
Xoutput160 net160 VGND VGND VPWR VPWR icache_adr_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput182 net182 VGND VGND VPWR VPWR store_data_o[23] sky130_fd_sc_hd__buf_4
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10070_ u_rf.reg9_q\[15\] _04459_ _04838_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__mux2_1
Xoutput171 net171 VGND VGND VPWR VPWR store_data_o[13] sky130_fd_sc_hd__clkbuf_4
Xoutput193 net193 VGND VGND VPWR VPWR store_data_o[4] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10972_ _05339_ VGND VGND VPWR VPWR _00709_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12711_ clknet_leaf_5_clk _00748_ net214 VGND VGND VPWR VPWR u_rf.reg23_q\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_48_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12642_ clknet_leaf_130_clk _00679_ net235 VGND VGND VPWR VPWR u_rf.reg21_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12573_ clknet_leaf_14_clk _00610_ net244 VGND VGND VPWR VPWR u_rf.reg19_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_525 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11524_ _05631_ VGND VGND VPWR VPWR _00969_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11455_ _04740_ u_rf.reg29_q\[9\] _05585_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10406_ _04782_ u_rf.reg13_q\[29\] _05028_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _05558_ VGND VGND VPWR VPWR _00904_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10337_ _05000_ VGND VGND VPWR VPWR _00413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10268_ u_rf.reg12_q\[7\] _04953_ _04939_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__mux2_1
X_12007_ clknet_leaf_79_clk u_exe.bu_pc_res\[20\] net372 VGND VGND VPWR VPWR u_exe.pc_data_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10199_ _04745_ u_rf.reg11_q\[11\] _04911_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12909_ clknet_leaf_8_clk _00946_ net226 VGND VGND VPWR VPWR u_rf.reg29_q\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06430_ u_decod.rs1_data_q\[1\] _01493_ _01428_ _01484_ u_decod.pc_q_o\[1\] VGND
+ VGND VPWR VPWR _01699_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06361_ _01630_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06292_ _01561_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__buf_8
X_08100_ _03235_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__buf_8
X_09080_ _04210_ _04217_ _04214_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__or3_1
XFILLER_0_72_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_96_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08031_ _03170_ _03209_ _03198_ VGND VGND VPWR VPWR _03237_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_79_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_761 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 load_data_i[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_142_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput73 reset_adr_i[17] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput62 load_data_i[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput51 load_data_i[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput84 reset_adr_i[27] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_0_141_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput95 reset_adr_i[8] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09982_ u_rf.reg8_q\[6\] _04440_ _04790_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08933_ _01380_ u_decod.branch_imm_q_o\[17\] VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__xor2_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08864_ _04030_ _04031_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__nor2_1
X_07815_ _03022_ _03024_ _03026_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_127_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ u_rf.reg30_q\[29\] _03280_ _03325_ u_rf.reg5_q\[29\] _03969_ VGND VGND VPWR
+ VPWR _03970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07746_ _02723_ _02922_ _02962_ _01443_ VGND VGND VPWR VPWR _02963_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_140_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09416_ u_decod.rf_ff_res_data_i\[21\] VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__buf_2
X_07677_ u_rf.reg18_q\[25\] _01592_ _01638_ u_rf.reg21_q\[25\] _02896_ VGND VGND VPWR
+ VPWR _02897_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06628_ u_rf.reg16_q\[4\] _01564_ _01630_ u_rf.reg17_q\[4\] VGND VGND VPWR VPWR _01890_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09347_ u_decod.rf_ff_rd_adr_q_i\[1\] VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_43_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06559_ _01444_ _01823_ _01497_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09278_ u_decod.instr_unit_q\[3\] VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__buf_2
XFILLER_0_132_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08229_ u_rf.reg1_q\[3\] _03311_ _03313_ u_rf.reg14_q\[3\] VGND VGND VPWR VPWR _03430_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11240_ _05481_ VGND VGND VPWR VPWR _00835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11171_ u_rf.reg25_q\[3\] _04945_ _05441_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__mux2_1
X_10122_ _04871_ VGND VGND VPWR VPWR _00327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10053_ u_rf.reg9_q\[7\] _04442_ _04827_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10955_ u_rf.reg21_q\[30\] _05001_ _05296_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10886_ u_rf.reg20_q\[30\] _05001_ _05259_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12625_ clknet_leaf_54_clk _00662_ net296 VGND VGND VPWR VPWR u_rf.reg20_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12556_ clknet_leaf_9_clk _00593_ net225 VGND VGND VPWR VPWR u_rf.reg18_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ _04724_ u_rf.reg30_q\[1\] _05621_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12487_ clknet_leaf_3_clk _00524_ net213 VGND VGND VPWR VPWR u_rf.reg16_q\[12\] sky130_fd_sc_hd__dfrtp_1
Xhold109 u_exe.pc_data_q\[11\] VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _05586_ VGND VGND VPWR VPWR _00928_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11369_ u_rf.reg28_q\[0\] net503 _05549_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_88 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05930_ _01216_ VGND VGND VPWR VPWR u_decod.dec0.rd_o\[2\] sky130_fd_sc_hd__clkbuf_1
X_05861_ u_decod.pc0_q_i\[20\] _01159_ VGND VGND VPWR VPWR _01163_ sky130_fd_sc_hd__or2_1
X_07600_ u_decod.rs2_data_q\[24\] u_decod.rs1_data_q\[24\] _02781_ VGND VGND VPWR
+ VPWR _02823_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08580_ u_rf.reg16_q\[19\] _03323_ _03325_ u_rf.reg5_q\[19\] _03764_ VGND VGND VPWR
+ VPWR _03765_ sky130_fd_sc_hd__a221o_1
X_07531_ u_rf.reg5_q\[22\] _02664_ _02375_ u_rf.reg11_q\[22\] _02756_ VGND VGND VPWR
+ VPWR _02757_ sky130_fd_sc_hd__a221o_1
X_05792_ u_decod.pc0_q_i\[2\] u_decod.pc0_q_i\[3\] u_decod.pc0_q_i\[4\] VGND VGND
+ VPWR VPWR _01110_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07462_ _02619_ net46 VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09201_ _04112_ _04274_ _04320_ _04322_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[20\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07393_ _02455_ _02623_ _01472_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__mux2_1
X_06413_ _01511_ _01528_ _01682_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[0\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09132_ u_decod.pc_q_o\[11\] u_decod.branch_imm_q_o\[11\] VGND VGND VPWR VPWR _04263_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06344_ _01538_ _01558_ _01577_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__and3_2
XFILLER_0_115_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09063_ _04202_ _04203_ VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__and2b_1
X_06275_ _01542_ u_decod.dec0.instr_i\[21\] _01544_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08014_ u_rf.reg22_q\[31\] _03218_ _03219_ u_rf.reg3_q\[31\] VGND VGND VPWR VPWR
+ _03220_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09965_ _04786_ u_rf.reg7_q\[31\] _04721_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08916_ _04062_ _04065_ _04069_ _04076_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a31o_1
X_09896_ u_decod.rf_ff_res_data_i\[9\] VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__buf_2
X_08847_ _03998_ _04017_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__nor2_1
X_08778_ _03944_ _03953_ _03378_ VGND VGND VPWR VPWR _03954_ sky130_fd_sc_hd__o21a_1
X_07729_ u_rf.reg25_q\[26\] _01783_ _02364_ u_rf.reg21_q\[26\] _02946_ VGND VGND VPWR
+ VPWR _02947_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ u_rf.reg18_q\[25\] _04991_ _05210_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10671_ _05179_ VGND VGND VPWR VPWR _00568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12410_ clknet_leaf_61_clk _00447_ net343 VGND VGND VPWR VPWR u_rf.reg13_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ clknet_leaf_46_clk _00378_ net298 VGND VGND VPWR VPWR u_rf.reg11_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12272_ clknet_leaf_34_clk _00309_ net275 VGND VGND VPWR VPWR u_rf.reg9_q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11223_ u_rf.reg25_q\[28\] _04997_ _05463_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ _05435_ VGND VGND VPWR VPWR _00795_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11085_ _04778_ u_rf.reg23_q\[27\] _05391_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__mux2_1
X_10105_ _04643_ _04682_ _04825_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__and3_4
X_10036_ _01531_ _01535_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11987_ clknet_leaf_88_clk u_exe.bu_pc_res\[0\] net360 VGND VGND VPWR VPWR u_exe.pc_data_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10938_ _05321_ VGND VGND VPWR VPWR _00693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10869_ _05284_ VGND VGND VPWR VPWR _00661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12608_ clknet_leaf_116_clk _00645_ net324 VGND VGND VPWR VPWR u_rf.reg20_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12539_ clknet_leaf_12_clk _00576_ net243 VGND VGND VPWR VPWR u_rf.reg18_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_563 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06060_ _01324_ _01327_ _01330_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__and3_1
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06962_ u_rf.reg1_q\[11\] _01587_ _01606_ u_rf.reg3_q\[11\] _02209_ VGND VGND VPWR
+ VPWR _02210_ sky130_fd_sc_hd__a221o_1
X_09750_ _04657_ VGND VGND VPWR VPWR _00169_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ u_rf.reg26_q\[25\] _03343_ _03285_ u_rf.reg21_q\[25\] VGND VGND VPWR VPWR
+ _03880_ sky130_fd_sc_hd__a22o_1
X_05913_ _01202_ VGND VGND VPWR VPWR _01203_ sky130_fd_sc_hd__inv_2
X_09681_ u_rf.reg4_q\[10\] _04448_ _04619_ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08632_ net443 _03773_ _03814_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[21\]
+ sky130_fd_sc_hd__a22o_1
X_06893_ _01458_ _02142_ _02143_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05844_ u_decod.pc0_q_i\[15\] u_decod.pc0_q_i\[16\] _01143_ VGND VGND VPWR VPWR _01150_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08563_ _03742_ _03744_ _03746_ _03748_ VGND VGND VPWR VPWR _03749_ sky130_fd_sc_hd__or4_1
X_05775_ _01097_ VGND VGND VPWR VPWR u_decod.dec0.unsign_extension sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08494_ u_rf.reg15_q\[15\] _03301_ _03303_ u_rf.reg24_q\[15\] _03682_ VGND VGND VPWR
+ VPWR _03683_ sky130_fd_sc_hd__a221o_1
X_07514_ _01437_ _02737_ _02738_ _02740_ VGND VGND VPWR VPWR _02741_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07445_ _01405_ _02635_ _01366_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_72 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07376_ u_rf.reg29_q\[19\] _01628_ _01659_ u_rf.reg14_q\[19\] _02607_ VGND VGND VPWR
+ VPWR _02608_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09115_ _04246_ _04248_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06327_ _01596_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__buf_8
XFILLER_0_33_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ u_decod.unsign_ext_q_o _04188_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__nand2_1
X_06258_ _01518_ _01527_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__or2_4
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06189_ _01444_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09948_ _04775_ VGND VGND VPWR VPWR _00249_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _04728_ u_rf.reg7_q\[3\] _04722_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__mux2_1
X_12890_ clknet_leaf_94_clk _00927_ net344 VGND VGND VPWR VPWR u_rf.reg28_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_11910_ clknet_leaf_91_clk u_decod.rs2_data_nxt\[31\] net345 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11841_ clknet_leaf_131_clk _00068_ net227 VGND VGND VPWR VPWR u_rf.reg0_q\[4\] sky130_fd_sc_hd__dfrtp_1
X_11772_ clknet_leaf_76_clk net369 net369 VGND VGND VPWR VPWR u_ifetch.reset_n_q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10723_ net519 _04974_ _05199_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10654_ _05170_ VGND VGND VPWR VPWR _00560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10585_ u_rf.reg16_q\[16\] _04972_ _05127_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_656 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12324_ clknet_leaf_109_clk _00361_ net313 VGND VGND VPWR VPWR u_rf.reg11_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12255_ clknet_leaf_131_clk _00292_ net227 VGND VGND VPWR VPWR u_rf.reg9_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11206_ _05440_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__buf_6
XFILLER_0_102_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12186_ clknet_leaf_61_clk _00223_ net341 VGND VGND VPWR VPWR u_rf.reg6_q\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _05426_ VGND VGND VPWR VPWR _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11068_ _04761_ u_rf.reg23_q\[19\] _05380_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__mux2_1
X_10019_ _04816_ VGND VGND VPWR VPWR _00279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_614 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07230_ u_rf.reg25_q\[16\] _01575_ _01624_ u_rf.reg28_q\[16\] VGND VGND VPWR VPWR
+ _02468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07161_ _02249_ _02295_ _02340_ _02401_ _02189_ _01476_ VGND VGND VPWR VPWR _02402_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06112_ _01381_ _01382_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07092_ u_decod.pc_q_o\[12\] u_decod.pc_q_o\[13\] u_decod.pc_q_o\[14\] _02185_ VGND
+ VGND VPWR VPWR _02335_ sky130_fd_sc_hd__and4_2
X_06043_ u_decod.rs1_data_q\[0\] u_decod.rs2_data_q\[0\] VGND VGND VPWR VPWR _01314_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout205 net206 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout216 net219 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_4
Xfanout238 net254 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_2
Xfanout227 net228 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_4
X_09802_ net522 _04430_ _04684_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07994_ _03188_ _03198_ _03199_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__and3_4
XFILLER_0_66_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout249 net252 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_105_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06945_ _02101_ _02193_ _01757_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__mux2_1
X_09733_ u_rf.reg5_q\[1\] _04430_ _04647_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_1
X_09664_ u_rf.reg4_q\[2\] _04432_ _04608_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__mux2_1
X_06876_ u_rf.reg1_q\[9\] _01585_ _01634_ u_rf.reg9_q\[9\] _02127_ VGND VGND VPWR
+ VPWR _02128_ sky130_fd_sc_hd__a221o_1
X_08615_ u_rf.reg18_q\[21\] _03353_ _03355_ u_rf.reg23_q\[21\] _03797_ VGND VGND VPWR
+ VPWR _03798_ sky130_fd_sc_hd__a221o_1
X_05827_ u_decod.pc0_q_i\[12\] _01133_ VGND VGND VPWR VPWR _01137_ sky130_fd_sc_hd__nand2_1
X_09595_ u_rf.reg3_q\[2\] _04432_ _04571_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__mux2_1
X_08546_ u_rf.reg6_q\[18\] _03304_ _03225_ u_rf.reg17_q\[18\] VGND VGND VPWR VPWR
+ _03732_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05758_ u_decod.dec0.funct7\[1\] u_decod.dec0.funct7\[0\] VGND VGND VPWR VPWR _01081_
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_137_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ u_decod.rf_ff_res_data_i\[14\] _03382_ _03666_ _03404_ VGND VGND VPWR VPWR
+ _03667_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_748 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07428_ u_rf.reg26_q\[20\] _01642_ _01645_ u_rf.reg20_q\[20\] VGND VGND VPWR VPWR
+ _02658_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_114_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07359_ _01443_ _02582_ _02591_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10370_ _05019_ VGND VGND VPWR VPWR _00427_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09029_ _01267_ u_decod.branch_imm_q_o\[31\] VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12040_ clknet_leaf_66_clk u_decod.exe_ff_res_data_i\[20\] net355 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[20\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_53_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_123_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ clknet_leaf_7_clk _00979_ net218 VGND VGND VPWR VPWR u_rf.reg30_q\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_143 _03265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net310 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ clknet_leaf_20_clk _00910_ net283 VGND VGND VPWR VPWR u_rf.reg28_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_132 _01625_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_110 u_decod.rs1_data_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11824_ clknet_leaf_93_clk net11 net344 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_165 u_decod.pc0_q_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 _03388_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_132_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11755_ clknet_leaf_29_clk _00047_ net257 VGND VGND VPWR VPWR u_rf.reg1_q\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_198 u_decod.rs1_data_q\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_187 _01605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ u_rf.reg18_q\[9\] _04957_ _05188_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11686_ u_decod.branch_imm_q_o\[21\] _02696_ _05717_ VGND VGND VPWR VPWR _05718_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10637_ _05161_ VGND VGND VPWR VPWR _00552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10568_ u_rf.reg16_q\[8\] _04955_ _05116_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__mux2_1
X_12307_ clknet_leaf_54_clk _00344_ net303 VGND VGND VPWR VPWR u_rf.reg10_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10499_ _05087_ VGND VGND VPWR VPWR _00488_ sky130_fd_sc_hd__clkbuf_1
X_12238_ clknet_leaf_28_clk _00275_ net256 VGND VGND VPWR VPWR u_rf.reg8_q\[19\] sky130_fd_sc_hd__dfrtp_1
X_12169_ clknet_leaf_24_clk _00206_ net267 VGND VGND VPWR VPWR u_rf.reg6_q\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06730_ u_decod.dec0.funct7\[1\] _01530_ _01548_ u_decod.rf_ff_res_data_i\[6\] VGND
+ VGND VPWR VPWR _01988_ sky130_fd_sc_hd__a22o_1
Xinput5 icache_instr_i[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_06661_ _01908_ _01913_ _01921_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08400_ u_rf.reg26_q\[11\] _03284_ _03345_ u_rf.reg21_q\[11\] VGND VGND VPWR VPWR
+ _03593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06592_ net36 _01489_ _01490_ net53 VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__a22o_1
X_09380_ _04447_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
X_08331_ u_rf.reg26_q\[8\] _03284_ _03286_ u_rf.reg21_q\[8\] VGND VGND VPWR VPWR _03527_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08262_ u_rf.reg6_q\[5\] _03387_ _03295_ u_rf.reg20_q\[5\] _03460_ VGND VGND VPWR
+ VPWR _03461_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07213_ _01763_ _02244_ _01400_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08193_ u_rf.reg30_q\[2\] _03280_ _03282_ u_rf.reg10_q\[2\] _03394_ VGND VGND VPWR
+ VPWR _03395_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07144_ _01671_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_399 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07075_ u_rf.reg23_q\[13\] _01612_ _01621_ u_rf.reg24_q\[13\] VGND VGND VPWR VPWR
+ _02319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06026_ u_decod.rs1_data_q\[12\] VGND VGND VPWR VPWR _01297_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07977_ _03180_ u_decod.exe_ff_rd_adr_q_i\[0\] u_decod.exe_ff_rd_adr_q_i\[4\] _03171_
+ _03182_ VGND VGND VPWR VPWR _03183_ sky130_fd_sc_hd__a221o_1
X_09716_ u_rf.reg4_q\[27\] _04484_ _04630_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__mux2_1
X_06928_ _02084_ _02132_ VGND VGND VPWR VPWR _02178_ sky130_fd_sc_hd__or2_1
X_09647_ u_rf.reg3_q\[27\] _04484_ _04593_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06859_ _02111_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[9\] sky130_fd_sc_hd__inv_2
X_09578_ _04563_ VGND VGND VPWR VPWR _00091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08529_ u_rf.reg18_q\[17\] _03352_ _03354_ u_rf.reg23_q\[17\] _03715_ VGND VGND VPWR
+ VPWR _03716_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11540_ _04757_ u_rf.reg30_q\[17\] _05632_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _05603_ VGND VGND VPWR VPWR _00944_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10422_ _04730_ u_rf.reg14_q\[4\] _05042_ VGND VGND VPWR VPWR _05047_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_458 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10353_ _05010_ VGND VGND VPWR VPWR _00419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10284_ u_rf.reg12_q\[12\] _04964_ _04960_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__mux2_1
X_12023_ clknet_leaf_114_clk u_decod.exe_ff_res_data_i\[3\] net328 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12925_ clknet_leaf_15_clk _00962_ net252 VGND VGND VPWR VPWR u_rf.reg30_q\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_53_clk _00893_ net304 VGND VGND VPWR VPWR u_rf.reg27_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11807_ clknet_leaf_106_clk net23 net320 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12787_ clknet_leaf_68_clk _00824_ net350 VGND VGND VPWR VPWR u_rf.reg25_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11738_ clknet_leaf_62_clk _00030_ net343 VGND VGND VPWR VPWR u_rf.reg2_q\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11669_ _05700_ net486 VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07900_ u_rf.reg0_q\[30\] _01664_ _01668_ u_rf.reg8_q\[30\] VGND VGND VPWR VPWR _03110_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_110_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08880_ _04037_ _04040_ _04036_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07831_ _01266_ _03003_ _01264_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__a21oi_1
X_09501_ _04522_ VGND VGND VPWR VPWR _00055_ sky130_fd_sc_hd__clkbuf_1
X_07762_ u_rf.reg6_q\[27\] _01557_ _02375_ u_rf.reg11_q\[27\] VGND VGND VPWR VPWR
+ _02978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07693_ _01357_ _01393_ _01407_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__a21o_1
X_06713_ u_rf.reg17_q\[6\] _01629_ _01652_ u_rf.reg22_q\[6\] VGND VGND VPWR VPWR _01971_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09432_ u_rf.reg2_q\[26\] _04482_ _04470_ VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__mux2_1
X_06644_ _01458_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09363_ u_decod.rf_ff_res_data_i\[4\] VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__buf_2
X_06575_ u_rf.reg15_q\[3\] _01600_ _01621_ u_rf.reg24_q\[3\] VGND VGND VPWR VPWR _01839_
+ sky130_fd_sc_hd__a22o_1
X_08314_ u_rf.reg6_q\[7\] _03305_ _03307_ u_rf.reg13_q\[7\] VGND VGND VPWR VPWR _03511_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_32 _03264_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _01597_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_21 _01679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09294_ _04385_ u_decod.rs2_data_q\[10\] _04386_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__and3_1
XANTENNA_65 _03428_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _03295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_54 _03337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08245_ u_rf.reg15_q\[4\] _03301_ _03303_ u_rf.reg24_q\[4\] _03444_ VGND VGND VPWR
+ VPWR _03445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_76 _04764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 _05585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _05152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08176_ _03347_ _03362_ _03377_ _03378_ VGND VGND VPWR VPWR _03379_ sky130_fd_sc_hd__o31a_1
X_07127_ u_rf.reg7_q\[14\] _01561_ _02368_ u_rf.reg26_q\[14\] VGND VGND VPWR VPWR
+ _02369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput150 net150 VGND VGND VPWR VPWR icache_adr_o[24] sky130_fd_sc_hd__buf_4
XFILLER_0_101_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput161 net161 VGND VGND VPWR VPWR icache_adr_o[5] sky130_fd_sc_hd__buf_2
X_07058_ _01441_ _02291_ _02298_ _02302_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__a211o_1
XFILLER_0_2_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput183 net183 VGND VGND VPWR VPWR store_data_o[24] sky130_fd_sc_hd__clkbuf_4
X_06009_ _01278_ _01279_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__and2_2
Xoutput172 net172 VGND VGND VPWR VPWR store_data_o[14] sky130_fd_sc_hd__clkbuf_4
Xoutput194 net194 VGND VGND VPWR VPWR store_data_o[5] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_145_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10971_ u_rf.reg22_q\[5\] _04949_ _05333_ VGND VGND VPWR VPWR _05339_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12710_ clknet_leaf_0_clk _00747_ net203 VGND VGND VPWR VPWR u_rf.reg23_q\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ clknet_leaf_95_clk _00678_ net327 VGND VGND VPWR VPWR u_rf.reg21_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ clknet_leaf_109_clk _00609_ net237 VGND VGND VPWR VPWR u_rf.reg19_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11523_ _04740_ u_rf.reg30_q\[9\] _05621_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__mux2_1
X_11454_ _05594_ VGND VGND VPWR VPWR _00936_ sky130_fd_sc_hd__clkbuf_1
X_10405_ _05037_ VGND VGND VPWR VPWR _00444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11385_ u_rf.reg28_q\[8\] u_decod.rf_ff_res_data_i\[8\] _05549_ VGND VGND VPWR VPWR
+ _05558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10336_ u_rf.reg12_q\[29\] _04999_ _04981_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10267_ u_decod.rf_ff_res_data_i\[7\] VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__buf_2
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_12006_ clknet_leaf_79_clk u_exe.bu_pc_res\[19\] net372 VGND VGND VPWR VPWR u_exe.pc_data_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10198_ _04912_ VGND VGND VPWR VPWR _00362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12908_ clknet_leaf_9_clk _00945_ net225 VGND VGND VPWR VPWR u_rf.reg29_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12839_ clknet_leaf_2_clk _00876_ net214 VGND VGND VPWR VPWR u_rf.reg27_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06360_ _01629_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06291_ _01560_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__buf_6
XFILLER_0_44_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08030_ _03171_ _03198_ _03204_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__and3_4
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput30 icache_instr_i[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_96_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput63 load_data_i[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
XFILLER_0_4_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput41 load_data_i[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput52 load_data_i[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_2
XFILLER_0_25_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput85 reset_adr_i[28] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XFILLER_0_141_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput74 reset_adr_i[18] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
Xinput96 reset_adr_i[9] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09981_ _04796_ VGND VGND VPWR VPWR _00261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08932_ _04042_ _04090_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08863_ u_decod.rs1_data_q\[7\] u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _04031_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_35_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07814_ u_rf.reg0_q\[28\] _01664_ _02371_ u_rf.reg15_q\[28\] _03027_ VGND VGND VPWR
+ VPWR _03028_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08794_ u_rf.reg16_q\[29\] _03322_ _03318_ u_rf.reg27_q\[29\] VGND VGND VPWR VPWR
+ _03969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07745_ _02723_ _02961_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_140_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ _04471_ VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__clkbuf_1
X_07676_ u_rf.reg25_q\[25\] _01575_ _01621_ u_rf.reg24_q\[25\] VGND VGND VPWR VPWR
+ _02896_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_180 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06627_ u_rf.reg0_q\[4\] _01662_ _01601_ u_rf.reg15_q\[4\] _01888_ VGND VGND VPWR
+ VPWR _01889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09346_ _04422_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__buf_6
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06558_ _01702_ u_decod.rs1_data_q\[3\] _01703_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09277_ _02685_ _03998_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__nor2_2
X_06489_ _01453_ _01755_ _01464_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08228_ _03315_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__buf_8
XFILLER_0_62_345 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08159_ _03351_ _03359_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11170_ _05444_ VGND VGND VPWR VPWR _00802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10121_ u_rf.reg10_q\[7\] _04442_ _04863_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__mux2_1
X_10052_ _04834_ VGND VGND VPWR VPWR _00294_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10954_ _05329_ VGND VGND VPWR VPWR _00701_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10885_ _05292_ VGND VGND VPWR VPWR _00669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12624_ clknet_leaf_34_clk _00661_ net275 VGND VGND VPWR VPWR u_rf.reg20_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12555_ clknet_leaf_135_clk _00592_ net209 VGND VGND VPWR VPWR u_rf.reg18_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11506_ _05622_ VGND VGND VPWR VPWR _00960_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12486_ clknet_leaf_140_clk _00523_ net203 VGND VGND VPWR VPWR u_rf.reg16_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11437_ _04719_ u_rf.reg29_q\[0\] _05585_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11368_ _05548_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10319_ _04988_ VGND VGND VPWR VPWR _00407_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11299_ _01531_ _01535_ _04568_ _05113_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__or4_4
X_05860_ u_decod.pc0_q_i\[20\] _01159_ VGND VGND VPWR VPWR _01162_ sky130_fd_sc_hd__and2_4
XFILLER_0_28_98 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05791_ net513 _01105_ _01101_ net90 _01109_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__a221o_2
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07530_ u_rf.reg27_q\[22\] _01671_ _01667_ u_rf.reg8_q\[22\] VGND VGND VPWR VPWR
+ _02756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07461_ _01506_ _02687_ _02689_ _01260_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09200_ _04319_ _04321_ _04196_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__a21boi_1
X_07392_ _01468_ _02237_ _01498_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__o21a_1
X_06412_ u_decod.dec0.instr_i\[20\] _01530_ _01550_ u_decod.rf_ff_res_data_i\[0\]
+ _01681_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_134_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09131_ u_decod.pc_q_o\[11\] u_decod.branch_imm_q_o\[11\] VGND VGND VPWR VPWR _04262_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06343_ _01612_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__buf_6
XFILLER_0_127_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09062_ u_decod.branch_imm_q_o\[1\] u_decod.pc_q_o\[1\] VGND VGND VPWR VPWR _04203_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06274_ u_decod.flush_v u_decod.rf_write_v_q_i VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08013_ _03170_ _03173_ _03209_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__and3_2
XFILLER_0_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09964_ u_decod.rf_ff_res_data_i\[31\] VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__buf_2
X_08915_ _01297_ u_decod.branch_imm_q_o\[12\] _04075_ _04068_ VGND VGND VPWR VPWR
+ _04076_ sky130_fd_sc_hd__a31o_1
X_09895_ _04739_ VGND VGND VPWR VPWR _00232_ sky130_fd_sc_hd__clkbuf_1
X_08846_ _04014_ net407 VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__xnor2_1
X_08777_ _03946_ _03948_ _03950_ _03952_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__or4_1
X_05989_ _01259_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ u_rf.reg18_q\[26\] _01787_ _01784_ u_rf.reg24_q\[26\] VGND VGND VPWR VPWR
+ _02946_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07659_ net100 net50 VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10670_ u_rf.reg17_q\[24\] _04989_ _05174_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09329_ _04413_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__buf_1
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12340_ clknet_leaf_22_clk _00377_ net268 VGND VGND VPWR VPWR u_rf.reg11_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12271_ clknet_leaf_44_clk _00308_ net275 VGND VGND VPWR VPWR u_rf.reg9_q\[20\] sky130_fd_sc_hd__dfrtp_1
X_11222_ _05471_ VGND VGND VPWR VPWR _00827_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11153_ u_rf.reg24_q\[27\] _04995_ _05427_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11084_ _05398_ VGND VGND VPWR VPWR _00762_ sky130_fd_sc_hd__clkbuf_1
X_10104_ _04861_ VGND VGND VPWR VPWR _00319_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10035_ _04824_ VGND VGND VPWR VPWR _00287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11986_ clknet_leaf_103_clk u_decod.dec0.unit_o\[3\] net335 VGND VGND VPWR VPWR u_decod.instr_unit_q\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_156_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10937_ u_rf.reg21_q\[21\] _04983_ _05319_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10868_ u_rf.reg20_q\[21\] _04983_ _05282_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__mux2_1
X_12607_ clknet_leaf_132_clk _00644_ net228 VGND VGND VPWR VPWR u_rf.reg20_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10799_ _05247_ VGND VGND VPWR VPWR _00628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12538_ clknet_leaf_59_clk _00575_ net289 VGND VGND VPWR VPWR u_rf.reg17_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12469_ clknet_leaf_47_clk _00506_ net300 VGND VGND VPWR VPWR u_rf.reg15_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06961_ u_rf.reg12_q\[11\] _01608_ _01642_ u_rf.reg26_q\[11\] VGND VGND VPWR VPWR
+ _02209_ sky130_fd_sc_hd__a22o_1
X_08700_ u_rf.reg8_q\[25\] _03271_ _03273_ u_rf.reg29_q\[25\] _03878_ VGND VGND VPWR
+ VPWR _03879_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ _04607_ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__buf_8
X_05912_ _01201_ _01080_ u_decod.dec0.instr_i\[4\] VGND VGND VPWR VPWR _01202_ sky130_fd_sc_hd__or3b_1
XFILLER_0_146_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ u_decod.exe_ff_res_data_i\[21\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[21\]
+ _03813_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__a221o_1
X_06892_ _01460_ _01955_ _01498_ _01450_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__o211a_1
X_05843_ _01099_ _01147_ _01148_ _01149_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__a31o_1
X_08562_ u_rf.reg23_q\[18\] _03354_ _03313_ u_rf.reg14_q\[18\] _03747_ VGND VGND VPWR
+ VPWR _03748_ sky130_fd_sc_hd__a221o_1
X_05774_ _01071_ _01075_ _01078_ _01084_ _01096_ VGND VGND VPWR VPWR _01097_ sky130_fd_sc_hd__a41o_1
XFILLER_0_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08493_ u_rf.reg6_q\[15\] _03387_ _03388_ u_rf.reg13_q\[15\] VGND VGND VPWR VPWR
+ _03682_ sky130_fd_sc_hd__a22o_1
X_07513_ _01398_ _01429_ _01432_ _01372_ _02739_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07444_ _02671_ _02673_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[20\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_84 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07375_ u_rf.reg15_q\[19\] _01600_ _01644_ u_rf.reg20_q\[19\] VGND VGND VPWR VPWR
+ _02607_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09114_ _04241_ _04236_ _04238_ _04239_ _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__o311a_1
X_06326_ _01513_ _01566_ _01577_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__and3_2
XFILLER_0_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06257_ _01257_ _01519_ _01524_ _01526_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__or4_4
X_09045_ _04177_ _04187_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06188_ _01453_ _01456_ _01458_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__mux2_1
X_09947_ _04774_ u_rf.reg7_q\[25\] _04764_ VGND VGND VPWR VPWR _04775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ u_decod.rf_ff_res_data_i\[3\] VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__clkbuf_4
X_08829_ u_decod.rs1_data_q\[2\] u_decod.branch_imm_q_o\[2\] VGND VGND VPWR VPWR _04002_
+ sky130_fd_sc_hd__and2_1
X_11840_ clknet_leaf_124_clk _00067_ net231 VGND VGND VPWR VPWR u_rf.reg0_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11771_ clknet_leaf_94_clk _00063_ net339 VGND VGND VPWR VPWR u_rf.reg1_q\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10722_ _05206_ VGND VGND VPWR VPWR _00592_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10653_ u_rf.reg17_q\[16\] _04972_ _05163_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10584_ _05133_ VGND VGND VPWR VPWR _00527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12323_ clknet_leaf_108_clk _00360_ net313 VGND VGND VPWR VPWR u_rf.reg11_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12254_ clknet_leaf_124_clk _00291_ net231 VGND VGND VPWR VPWR u_rf.reg9_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_12185_ clknet_leaf_56_clk _00222_ net291 VGND VGND VPWR VPWR u_rf.reg6_q\[30\] sky130_fd_sc_hd__dfrtp_1
X_11205_ _05462_ VGND VGND VPWR VPWR _00819_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ u_rf.reg24_q\[19\] _04978_ _05416_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__mux2_1
X_11067_ _05389_ VGND VGND VPWR VPWR _00754_ sky130_fd_sc_hd__clkbuf_1
X_10018_ u_rf.reg8_q\[23\] _04476_ _04812_ VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11969_ clknet_leaf_79_clk net469 net372 VGND VGND VPWR VPWR u_decod.pc_q_o\[18\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_137_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_137_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_626 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_339 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07160_ _02197_ _02400_ _01905_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07091_ _01764_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__clkbuf_4
X_06111_ u_decod.rs2_data_q\[17\] _01380_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06042_ u_decod.rs1_data_q\[2\] u_decod.rs2_data_q\[2\] VGND VGND VPWR VPWR _01313_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09801_ _04685_ VGND VGND VPWR VPWR _00192_ sky130_fd_sc_hd__clkbuf_1
Xfanout217 net219 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout206 net207 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_2
Xfanout228 net233 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07993_ u_decod.dec0.instr_i\[15\] _03190_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__nor2_2
X_09732_ _04648_ VGND VGND VPWR VPWR _00160_ sky130_fd_sc_hd__clkbuf_1
Xfanout239 net254 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06944_ _01994_ _02192_ _01451_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__mux2_1
X_09663_ _04610_ VGND VGND VPWR VPWR _00129_ sky130_fd_sc_hd__clkbuf_1
X_06875_ u_rf.reg11_q\[9\] _01582_ _01665_ u_rf.reg8_q\[9\] VGND VGND VPWR VPWR _02127_
+ sky130_fd_sc_hd__a22o_1
X_08614_ u_rf.reg4_q\[21\] _03265_ _03267_ u_rf.reg17_q\[21\] VGND VGND VPWR VPWR
+ _03797_ sky130_fd_sc_hd__a22o_1
X_05826_ u_decod.pc0_q_i\[12\] _01133_ VGND VGND VPWR VPWR _01136_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09594_ _04573_ VGND VGND VPWR VPWR _00097_ sky130_fd_sc_hd__clkbuf_1
X_08545_ u_decod.pc0_q_i\[17\] _03565_ _03731_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[17\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_128_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_128_clk sky130_fd_sc_hd__clkbuf_16
X_05757_ u_decod.dec0.instr_i\[6\] VGND VGND VPWR VPWR _01080_ sky130_fd_sc_hd__buf_2
XFILLER_0_38_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08476_ _03649_ _03656_ _03665_ VGND VGND VPWR VPWR _03666_ sky130_fd_sc_hd__or3_2
XFILLER_0_64_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07427_ _02649_ _02651_ _02654_ _02656_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__or4_1
XFILLER_0_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07358_ _01059_ _02583_ _02587_ _02590_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06309_ _01578_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_150_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07289_ u_rf.reg29_q\[17\] _01627_ _01652_ u_rf.reg22_q\[17\] VGND VGND VPWR VPWR
+ _02525_ sky130_fd_sc_hd__a22o_1
X_09028_ _04168_ _04169_ _04166_ VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12941_ clknet_leaf_7_clk _00978_ net226 VGND VGND VPWR VPWR u_rf.reg30_q\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ clknet_leaf_17_clk _00909_ net288 VGND VGND VPWR VPWR u_rf.reg28_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_100 _05621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 u_decod.rs1_data_q\[26\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11823_ clknet_leaf_93_clk net10 net344 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_122 net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 _01656_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_155 _04695_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 u_decod.pc0_q_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_119_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_119_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_144 _03283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11754_ clknet_leaf_25_clk _00046_ net265 VGND VGND VPWR VPWR u_rf.reg1_q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_177 net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11685_ net357 VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_81_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10705_ _05197_ VGND VGND VPWR VPWR _00584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10636_ u_rf.reg17_q\[8\] _04955_ _05152_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10567_ _05124_ VGND VGND VPWR VPWR _00519_ sky130_fd_sc_hd__clkbuf_1
X_12306_ clknet_leaf_40_clk _00343_ net278 VGND VGND VPWR VPWR u_rf.reg10_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10498_ _04738_ u_rf.reg15_q\[8\] _05078_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12237_ clknet_leaf_6_clk _00274_ net215 VGND VGND VPWR VPWR u_rf.reg8_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ clknet_leaf_19_clk _00205_ net288 VGND VGND VPWR VPWR u_rf.reg6_q\[13\] sky130_fd_sc_hd__dfrtp_1
X_12099_ clknet_leaf_107_clk _00136_ net314 VGND VGND VPWR VPWR u_rf.reg4_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11119_ _05417_ VGND VGND VPWR VPWR _00778_ sky130_fd_sc_hd__clkbuf_1
Xinput6 icache_instr_i[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_06660_ _01310_ _01763_ _01916_ _01919_ _01920_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_149_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06591_ _01853_ _01854_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[3\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08330_ u_rf.reg8_q\[8\] _03271_ _03273_ u_rf.reg29_q\[8\] _03525_ VGND VGND VPWR
+ VPWR _03526_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08261_ u_rf.reg9_q\[5\] _03293_ _03216_ u_rf.reg8_q\[5\] VGND VGND VPWR VPWR _03460_
+ sky130_fd_sc_hd__a22o_1
X_07212_ _02295_ _02340_ _02401_ _02450_ _01478_ _01475_ VGND VGND VPWR VPWR _02451_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_15_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08192_ u_rf.reg26_q\[2\] _03203_ _03206_ u_rf.reg21_q\[2\] VGND VGND VPWR VPWR _03394_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07143_ _01645_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_132_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07074_ _02311_ _02313_ _02315_ _02317_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06025_ u_decod.rs2_data_q\[13\] u_decod.rs1_data_q\[13\] VGND VGND VPWR VPWR _01296_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07976_ u_decod.dec0.instr_i\[16\] _01521_ u_decod.exe_ff_rd_adr_q_i\[2\] _03181_
+ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__a22o_1
X_09715_ _04637_ VGND VGND VPWR VPWR _00154_ sky130_fd_sc_hd__clkbuf_1
X_06927_ _01713_ u_decod.exe_ff_res_data_i\[10\] _02176_ VGND VGND VPWR VPWR _02177_
+ sky130_fd_sc_hd__a21o_1
X_09646_ _04600_ VGND VGND VPWR VPWR _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_82 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06858_ _01765_ _02092_ _02097_ _02104_ _02110_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__o2111a_1
X_09577_ u_rf.reg0_q\[27\] _04484_ _04555_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__mux2_1
X_05809_ net478 _01105_ _01101_ net94 _01123_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__a221o_1
X_06789_ _01865_ _02043_ _01457_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__mux2_1
X_08528_ u_rf.reg4_q\[17\] _03264_ _03266_ u_rf.reg17_q\[17\] VGND VGND VPWR VPWR
+ _03715_ sky130_fd_sc_hd__a22o_1
X_08459_ u_rf.reg30_q\[14\] _03341_ _03342_ u_rf.reg10_q\[14\] _03648_ VGND VGND VPWR
+ VPWR _03649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11470_ _04755_ u_rf.reg29_q\[16\] _05596_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10421_ _05046_ VGND VGND VPWR VPWR _00451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10352_ _04728_ u_rf.reg13_q\[3\] _05006_ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12022_ clknet_leaf_97_clk u_decod.exe_ff_res_data_i\[2\] net331 VGND VGND VPWR VPWR
+ u_decod.rf_ff_res_data_i\[2\] sky130_fd_sc_hd__dfrtp_4
X_10283_ u_decod.rf_ff_res_data_i\[12\] VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_616 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12924_ clknet_leaf_126_clk _00961_ net240 VGND VGND VPWR VPWR u_rf.reg30_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ clknet_leaf_70_clk _00892_ net354 VGND VGND VPWR VPWR u_rf.reg27_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_12786_ clknet_leaf_38_clk _00823_ net274 VGND VGND VPWR VPWR u_rf.reg25_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11806_ clknet_leaf_106_clk net12 net320 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11737_ clknet_leaf_67_clk _00029_ net355 VGND VGND VPWR VPWR u_rf.reg2_q\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11668_ _05708_ VGND VGND VPWR VPWR _01036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10619_ _05151_ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__buf_6
XFILLER_0_52_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11599_ _05671_ VGND VGND VPWR VPWR _01004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07830_ _03041_ _03043_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[28\] sky130_fd_sc_hd__xnor2_1
X_07761_ u_rf.reg12_q\[27\] _01610_ _02697_ u_rf.reg4_q\[27\] _02976_ VGND VGND VPWR
+ VPWR _02977_ sky130_fd_sc_hd__a221o_1
X_09500_ net526 _04476_ _04518_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06712_ u_rf.reg11_q\[6\] _01583_ _01656_ u_rf.reg10_q\[6\] _01969_ VGND VGND VPWR
+ VPWR _01970_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07692_ _01276_ _01278_ _02821_ _02910_ _01410_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__a311o_1
XFILLER_0_63_30 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09431_ u_decod.rf_ff_res_data_i\[26\] VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06643_ _01444_ _01903_ _01497_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__o21a_1
X_06574_ u_rf.reg29_q\[3\] _01628_ _01667_ u_rf.reg8_q\[3\] _01837_ VGND VGND VPWR
+ VPWR _01838_ sky130_fd_sc_hd__a221o_1
X_09362_ _04435_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08313_ _03501_ _03503_ _03507_ _03509_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_11 _01600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09293_ _04393_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_1
XANTENNA_22 _01679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_44 _03295_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _03265_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _03343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 _03429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08244_ u_rf.reg6_q\[4\] _03305_ _03307_ u_rf.reg13_q\[4\] VGND VGND VPWR VPWR _03444_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_77 _04764_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _05246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08175_ _03253_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__buf_6
XANTENNA_99 _05585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07126_ _01642_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput151 net151 VGND VGND VPWR VPWR icache_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput140 net140 VGND VGND VPWR VPWR icache_adr_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_112_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07057_ _01295_ _01429_ _02299_ _01058_ _02301_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__a221o_1
Xoutput184 net184 VGND VGND VPWR VPWR store_data_o[25] sky130_fd_sc_hd__clkbuf_4
X_06008_ u_decod.rs2_data_q\[24\] u_decod.rs1_data_q\[24\] VGND VGND VPWR VPWR _01279_
+ sky130_fd_sc_hd__or2_1
Xoutput173 net173 VGND VGND VPWR VPWR store_data_o[15] sky130_fd_sc_hd__clkbuf_4
Xoutput195 net195 VGND VGND VPWR VPWR store_data_o[6] sky130_fd_sc_hd__clkbuf_4
Xoutput162 net162 VGND VGND VPWR VPWR icache_adr_o[6] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_145_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07959_ u_decod.dec0.unsign_extension _02229_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10970_ _05338_ VGND VGND VPWR VPWR _00708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09629_ _04591_ VGND VGND VPWR VPWR _00114_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ clknet_leaf_119_clk _00677_ net248 VGND VGND VPWR VPWR u_rf.reg21_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ clknet_leaf_11_clk _00608_ net222 VGND VGND VPWR VPWR u_rf.reg19_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11522_ _05630_ VGND VGND VPWR VPWR _00968_ sky130_fd_sc_hd__clkbuf_1
X_11453_ _04738_ u_rf.reg29_q\[8\] _05585_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10404_ _04780_ u_rf.reg13_q\[28\] _05028_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11384_ _05557_ VGND VGND VPWR VPWR _00903_ sky130_fd_sc_hd__clkbuf_1
X_10335_ u_decod.rf_ff_res_data_i\[29\] VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__buf_2
XFILLER_0_104_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10266_ _04952_ VGND VGND VPWR VPWR _00390_ sky130_fd_sc_hd__clkbuf_1
X_12005_ clknet_leaf_83_clk u_exe.bu_pc_res\[18\] net370 VGND VGND VPWR VPWR u_exe.pc_data_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10197_ _04742_ u_rf.reg11_q\[10\] _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12907_ clknet_leaf_1_clk _00944_ net209 VGND VGND VPWR VPWR u_rf.reg29_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12838_ clknet_leaf_0_clk _00875_ net204 VGND VGND VPWR VPWR u_rf.reg27_q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_546 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12769_ clknet_leaf_119_clk _00806_ net251 VGND VGND VPWR VPWR u_rf.reg25_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06290_ _01559_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__buf_8
XFILLER_0_154_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput31 icache_instr_i[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_4_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 icache_instr_i[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
XFILLER_0_142_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput64 load_data_i[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 load_data_i[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
XFILLER_0_4_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 load_data_i[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput75 reset_adr_i[19] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
Xinput86 reset_adr_i[29] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput97 reset_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
XFILLER_0_40_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09980_ u_rf.reg8_q\[5\] _04438_ _04790_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08931_ _04086_ net378 VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08862_ u_decod.rs1_data_q\[7\] u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _04030_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07813_ u_rf.reg30_q\[28\] _01581_ _02419_ u_rf.reg28_q\[28\] VGND VGND VPWR VPWR
+ _03027_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_150_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08793_ u_rf.reg8_q\[29\] _03270_ _03272_ u_rf.reg29_q\[29\] _03967_ VGND VGND VPWR
+ VPWR _03968_ sky130_fd_sc_hd__a221o_1
X_07744_ _02871_ _02960_ _02681_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07675_ u_rf.reg31_q\[25\] _01616_ _01658_ u_rf.reg14_q\[25\] _02894_ VGND VGND VPWR
+ VPWR _02895_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_140_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09414_ u_rf.reg2_q\[20\] _04469_ _04470_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06626_ u_rf.reg7_q\[4\] _01560_ _01605_ u_rf.reg3_q\[4\] VGND VGND VPWR VPWR _01888_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
X_09345_ _01539_ u_decod.rf_write_v_q_i VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06557_ _01815_ _01818_ _01821_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__or3b_1
X_09276_ _01477_ _03998_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__nor2_2
XFILLER_0_75_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06488_ _01752_ _01754_ _01467_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08227_ _03314_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__buf_8
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08158_ u_rf.reg8_q\[1\] _03271_ _03273_ u_rf.reg29_q\[1\] _03360_ VGND VGND VPWR
+ VPWR _03361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08089_ _03212_ VGND VGND VPWR VPWR _03293_ sky130_fd_sc_hd__buf_6
X_07109_ _01425_ _02351_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10120_ _04870_ VGND VGND VPWR VPWR _00326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10051_ u_rf.reg9_q\[6\] _04440_ _04827_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_99_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10953_ u_rf.reg21_q\[29\] _04999_ _05319_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10884_ u_rf.reg20_q\[29\] _04999_ _05282_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12623_ clknet_leaf_42_clk _00660_ net275 VGND VGND VPWR VPWR u_rf.reg20_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_23_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12554_ clknet_leaf_30_clk _00591_ net261 VGND VGND VPWR VPWR u_rf.reg18_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11505_ _04719_ u_rf.reg30_q\[0\] _05621_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ clknet_leaf_124_clk _00522_ net239 VGND VGND VPWR VPWR u_rf.reg16_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11436_ _05584_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11367_ _04937_ _05114_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__nor2_4
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10318_ u_rf.reg12_q\[23\] _04987_ _04981_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11298_ _05511_ VGND VGND VPWR VPWR _00863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10249_ u_decod.rf_ff_res_data_i\[1\] VGND VGND VPWR VPWR _04941_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_109_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05790_ net390 u_decod.pc0_q_i\[3\] _01108_ VGND VGND VPWR VPWR _01109_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_122_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07460_ _01430_ _01360_ _01361_ u_decod.instr_operation_q\[3\] _02688_ VGND VGND
+ VPWR VPWR _02689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07391_ _02618_ _02620_ _02621_ VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__a21oi_1
X_06411_ _01619_ _01677_ _01680_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__o21a_2
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09130_ _04054_ _04207_ _04208_ _04261_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[10\]
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06342_ _01611_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__buf_12
XFILLER_0_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09061_ u_decod.branch_imm_q_o\[1\] u_decod.pc_q_o\[1\] VGND VGND VPWR VPWR _04202_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08012_ u_decod.dec0.instr_i\[19\] _03199_ _03205_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__and3_2
X_06273_ _01542_ u_decod.dec0.instr_i\[21\] _01512_ u_decod.rf_ff_rd_adr_q_i\[4\]
+ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09963_ _04785_ VGND VGND VPWR VPWR _00254_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08914_ u_decod.rs1_data_q\[13\] u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR
+ _04075_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09894_ _04738_ u_rf.reg7_q\[8\] _04722_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__mux2_1
X_08845_ _04008_ _04005_ _04009_ _04015_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__a31o_1
X_08776_ u_rf.reg0_q\[28\] _03420_ _03421_ u_rf.reg12_q\[28\] _03951_ VGND VGND VPWR
+ VPWR _03952_ sky130_fd_sc_hd__a221o_1
X_07727_ u_rf.reg31_q\[26\] _01777_ _02367_ u_rf.reg14_q\[26\] _02944_ VGND VGND VPWR
+ VPWR _02945_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_243 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05988_ _01258_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07658_ _01506_ _02876_ _02878_ _01260_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_67_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07589_ _02357_ u_decod.exe_ff_res_data_i\[23\] _02812_ VGND VGND VPWR VPWR _02813_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
X_06609_ _01506_ _01867_ _01871_ _01442_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__a22o_1
X_09328_ _04409_ u_decod.rs2_data_q\[25\] _04410_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09259_ u_decod.pc_q_o\[29\] u_decod.branch_imm_q_o\[29\] VGND VGND VPWR VPWR _04372_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12270_ clknet_leaf_28_clk _00307_ net256 VGND VGND VPWR VPWR u_rf.reg9_q\[19\] sky130_fd_sc_hd__dfrtp_1
X_11221_ u_rf.reg25_q\[27\] _04995_ _05463_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11152_ _05434_ VGND VGND VPWR VPWR _00794_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10103_ u_rf.reg9_q\[31\] _04492_ _04826_ VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11083_ _04776_ u_rf.reg23_q\[26\] _05391_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10034_ u_rf.reg8_q\[31\] _04492_ _04789_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11985_ clknet_leaf_103_clk u_decod.dec0.is_branch net336 VGND VGND VPWR VPWR u_decod.instr_unit_q\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10936_ _05320_ VGND VGND VPWR VPWR _00692_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10867_ _05283_ VGND VGND VPWR VPWR _00660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12606_ clknet_leaf_124_clk _00643_ net231 VGND VGND VPWR VPWR u_rf.reg20_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10798_ u_rf.reg19_q\[20\] _04980_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__mux2_1
X_12537_ clknet_leaf_56_clk _00574_ net293 VGND VGND VPWR VPWR u_rf.reg17_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12468_ clknet_leaf_31_clk _00505_ net261 VGND VGND VPWR VPWR u_rf.reg15_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11419_ u_rf.reg28_q\[24\] net477 _05571_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__mux2_1
X_12399_ clknet_leaf_36_clk _00436_ net273 VGND VGND VPWR VPWR u_rf.reg13_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_06960_ u_rf.reg28_q\[11\] _01625_ _01653_ u_rf.reg22_q\[11\] _02207_ VGND VGND VPWR
+ VPWR _02208_ sky130_fd_sc_hd__a221o_1
X_06891_ _01748_ _02141_ _01685_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__mux2_1
X_05911_ u_decod.dec0.instr_i\[0\] _01074_ VGND VGND VPWR VPWR _01201_ sky130_fd_sc_hd__nand2_1
X_08630_ _03803_ _03812_ _03378_ VGND VGND VPWR VPWR _03813_ sky130_fd_sc_hd__o21a_2
X_05842_ u_exe.pc_data_q\[15\] _01118_ _01119_ net71 VGND VGND VPWR VPWR _01149_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08561_ u_rf.reg0_q\[18\] _03174_ _03276_ u_rf.reg3_q\[18\] VGND VGND VPWR VPWR _03747_
+ sky130_fd_sc_hd__a22o_1
X_05773_ _01071_ _01089_ _01090_ _01091_ _01095_ VGND VGND VPWR VPWR _01096_ sky130_fd_sc_hd__a221o_1
X_07512_ _01374_ _02244_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nor2_1
X_08492_ u_rf.reg7_q\[15\] _03369_ _03370_ u_rf.reg25_q\[15\] _03680_ VGND VGND VPWR
+ VPWR _03681_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07443_ _02089_ _02487_ _02672_ net199 VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07374_ u_rf.reg1_q\[19\] _02604_ _01576_ u_rf.reg25_q\[19\] _02605_ VGND VGND VPWR
+ VPWR _02606_ sky130_fd_sc_hd__a221o_1
X_09113_ _04238_ u_decod.branch_imm_q_o\[6\] u_decod.pc_q_o\[6\] VGND VGND VPWR VPWR
+ _04247_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06325_ _01594_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06256_ u_decod.dec0.instr_i\[21\] _01521_ u_decod.exe_ff_rd_adr_q_i\[4\] _01513_
+ _01525_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__o221ai_2
X_09044_ _01324_ _04178_ _04185_ _04186_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__or4b_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06187_ _01457_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09946_ u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _04727_ VGND VGND VPWR VPWR _00226_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_51_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ u_decod.rs1_data_q\[2\] u_decod.branch_imm_q_o\[2\] VGND VGND VPWR VPWR _04001_
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08759_ net452 _03773_ _03935_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[27\]
+ sky130_fd_sc_hd__a22o_1
X_11770_ clknet_leaf_61_clk _00062_ net341 VGND VGND VPWR VPWR u_rf.reg1_q\[30\] sky130_fd_sc_hd__dfrtp_1
X_10721_ u_rf.reg18_q\[16\] _04972_ _05199_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10652_ _05169_ VGND VGND VPWR VPWR _00559_ sky130_fd_sc_hd__clkbuf_1
X_10583_ u_rf.reg16_q\[15\] _04970_ _05127_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ clknet_leaf_128_clk _00359_ net234 VGND VGND VPWR VPWR u_rf.reg11_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12253_ clknet_leaf_122_clk _00290_ net248 VGND VGND VPWR VPWR u_rf.reg9_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11204_ u_rf.reg25_q\[19\] _04978_ _05452_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__mux2_1
X_12184_ clknet_leaf_53_clk _00221_ net304 VGND VGND VPWR VPWR u_rf.reg6_q\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11135_ _05425_ VGND VGND VPWR VPWR _00786_ sky130_fd_sc_hd__clkbuf_1
X_11066_ _04759_ u_rf.reg23_q\[18\] _05380_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__mux2_1
X_10017_ _04815_ VGND VGND VPWR VPWR _00278_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_511 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ clknet_leaf_83_clk net461 net365 VGND VGND VPWR VPWR u_decod.pc_q_o\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11899_ clknet_leaf_91_clk u_decod.rs2_data_nxt\[20\] net345 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10919_ _05311_ VGND VGND VPWR VPWR _00684_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_912 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07090_ _02331_ _02332_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06110_ u_decod.rs2_data_q\[17\] _01380_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06041_ u_decod.rs1_data_q\[3\] u_decod.rs2_data_q\[3\] VGND VGND VPWR VPWR _01312_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07992_ _03181_ _03191_ VGND VGND VPWR VPWR _03198_ sky130_fd_sc_hd__nor2_2
Xfanout218 net219 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_2
X_09800_ u_rf.reg6_q\[0\] _04421_ _04684_ VGND VGND VPWR VPWR _04685_ sky130_fd_sc_hd__mux2_1
Xfanout207 net210 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_2
Xfanout229 net233 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_4
X_09731_ u_rf.reg5_q\[0\] _04421_ _04647_ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__mux2_1
X_06943_ _02190_ _02191_ _01455_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09662_ u_rf.reg4_q\[1\] _04430_ _04608_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__mux2_1
X_06874_ u_rf.reg23_q\[9\] _01611_ _01655_ u_rf.reg10_q\[9\] _02125_ VGND VGND VPWR
+ VPWR _02126_ sky130_fd_sc_hd__a221o_1
X_08613_ u_rf.reg8_q\[21\] _03407_ _03408_ u_rf.reg29_q\[21\] _03795_ VGND VGND VPWR
+ VPWR _03796_ sky130_fd_sc_hd__a221o_1
X_05825_ net483 _01105_ _01132_ net67 _01135_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__a221o_1
X_09593_ u_rf.reg3_q\[1\] _04430_ _04571_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08544_ u_decod.exe_ff_res_data_i\[17\] _03381_ _03730_ VGND VGND VPWR VPWR _03731_
+ sky130_fd_sc_hd__a21o_1
X_05756_ u_decod.dec0.funct7\[5\] VGND VGND VPWR VPWR _01079_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08475_ _03658_ _03660_ _03662_ _03664_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__or4_1
XFILLER_0_92_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ u_rf.reg9_q\[20\] _01636_ _01668_ u_rf.reg8_q\[20\] _02655_ VGND VGND VPWR
+ VPWR _02656_ sky130_fd_sc_hd__a221o_1
XFILLER_0_119_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07357_ u_decod.rs2_data_q\[19\] _01376_ _01429_ _02589_ VGND VGND VPWR VPWR _02590_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_33_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06308_ _01538_ _01553_ _01577_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_150_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09027_ _04171_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_115_373 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07288_ u_rf.reg11_q\[17\] _01583_ _01598_ u_rf.reg13_q\[17\] _02523_ VGND VGND VPWR
+ VPWR _02524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_28_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06239_ _01443_ _01482_ _01509_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09929_ _04762_ VGND VGND VPWR VPWR _00243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12940_ clknet_leaf_10_clk _00977_ net224 VGND VGND VPWR VPWR u_rf.reg30_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12871_ clknet_leaf_2_clk _00908_ net223 VGND VGND VPWR VPWR u_rf.reg28_q\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_29_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 _05632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ clknet_leaf_93_clk net9 net344 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[17\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_134 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 u_decod.rs1_data_q\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 _03292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 _04874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_167 u_decod.pc_q_o\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11753_ clknet_leaf_18_clk _00045_ net288 VGND VGND VPWR VPWR u_rf.reg1_q\[13\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_178 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_189 _01658_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11684_ _05716_ VGND VGND VPWR VPWR _01044_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ u_rf.reg18_q\[8\] _04955_ _05188_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10635_ _05160_ VGND VGND VPWR VPWR _00551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12305_ clknet_leaf_56_clk _00342_ net286 VGND VGND VPWR VPWR u_rf.reg10_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10566_ u_rf.reg16_q\[7\] _04953_ _05116_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10497_ _05086_ VGND VGND VPWR VPWR _00487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12236_ clknet_leaf_25_clk _00273_ net265 VGND VGND VPWR VPWR u_rf.reg8_q\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12167_ clknet_leaf_4_clk _00204_ net211 VGND VGND VPWR VPWR u_rf.reg6_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_11118_ u_rf.reg24_q\[10\] _04959_ _05416_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__mux2_1
X_12098_ clknet_leaf_131_clk _00135_ net229 VGND VGND VPWR VPWR u_rf.reg4_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11049_ _05368_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__buf_8
Xinput7 icache_instr_i[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06590_ _01802_ _01805_ _01744_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_143_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08260_ u_rf.reg15_q\[5\] _03300_ _03388_ u_rf.reg13_q\[5\] _03458_ VGND VGND VPWR
+ VPWR _03459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08191_ _03386_ _03390_ _03392_ VGND VGND VPWR VPWR _03393_ sky130_fd_sc_hd__or3_1
X_07211_ _02248_ _02449_ _01458_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07142_ u_rf.reg16_q\[14\] _02307_ _01776_ u_rf.reg2_q\[14\] _02383_ VGND VGND VPWR
+ VPWR _02384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07073_ u_rf.reg3_q\[13\] _01606_ _01639_ u_rf.reg21_q\[13\] _02316_ VGND VGND VPWR
+ VPWR _02317_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06024_ u_decod.rs2_data_q\[13\] u_decod.rs1_data_q\[13\] VGND VGND VPWR VPWR _01295_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_11_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07975_ u_decod.dec0.instr_i\[17\] VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__inv_2
X_09714_ u_rf.reg4_q\[26\] _04482_ _04630_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__mux2_1
X_06926_ u_decod.dec0.funct7\[5\] _01530_ _01548_ u_decod.rf_ff_res_data_i\[10\] _02175_
+ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__a221o_1
X_09645_ u_rf.reg3_q\[26\] _04482_ _04593_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06857_ _01057_ _02105_ _02107_ _02109_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__o211a_1
X_05808_ _01121_ _01106_ _01122_ VGND VGND VPWR VPWR _01123_ sky130_fd_sc_hd__and3b_1
XFILLER_0_93_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_143_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _04562_ VGND VGND VPWR VPWR _00090_ sky130_fd_sc_hd__clkbuf_1
X_06788_ _01495_ _02042_ _01684_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__mux2_1
X_08527_ u_rf.reg9_q\[17\] _03348_ _03349_ u_rf.reg20_q\[17\] _03713_ VGND VGND VPWR
+ VPWR _03714_ sky130_fd_sc_hd__a221o_1
X_05739_ _01064_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__inv_2
XFILLER_0_136_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_605 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08458_ u_rf.reg26_q\[14\] _03344_ _03345_ u_rf.reg21_q\[14\] VGND VGND VPWR VPWR
+ _03648_ sky130_fd_sc_hd__a22o_1
X_07409_ _01764_ _02638_ _02639_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_46_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_468 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08389_ _03576_ _03578_ _03580_ _03582_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__or4_1
X_10420_ _04728_ u_rf.reg14_q\[3\] _05042_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10351_ _05009_ VGND VGND VPWR VPWR _00418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10282_ _04963_ VGND VGND VPWR VPWR _00395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12021_ clknet_leaf_113_clk u_decod.exe_ff_res_data_i\[1\] net328 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[1\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_45_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12923_ clknet_leaf_13_clk _00960_ net242 VGND VGND VPWR VPWR u_rf.reg30_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12854_ clknet_leaf_48_clk _00891_ net306 VGND VGND VPWR VPWR u_rf.reg27_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12785_ clknet_leaf_56_clk _00822_ net287 VGND VGND VPWR VPWR u_rf.reg25_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11805_ clknet_leaf_105_clk net1 net320 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_11736_ clknet_leaf_72_clk _00028_ net353 VGND VGND VPWR VPWR u_rf.reg2_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11667_ u_decod.branch_imm_q_o\[12\] _02257_ _05696_ VGND VGND VPWR VPWR _05708_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10618_ _04494_ _05114_ VGND VGND VPWR VPWR _05151_ sky130_fd_sc_hd__nor2_4
X_11598_ _04747_ u_rf.reg31_q\[12\] _05668_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10549_ _05113_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__buf_6
XFILLER_0_51_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_63_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12219_ clknet_leaf_12_clk _00256_ net243 VGND VGND VPWR VPWR u_rf.reg8_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07760_ u_rf.reg31_q\[27\] _01777_ _02380_ u_rf.reg10_q\[27\] VGND VGND VPWR VPWR
+ _02976_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06711_ u_rf.reg9_q\[6\] _01635_ _01666_ u_rf.reg8_q\[6\] VGND VGND VPWR VPWR _01969_
+ sky130_fd_sc_hd__a22o_1
X_09430_ _04481_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__clkbuf_1
X_07691_ _01286_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06642_ u_decod.rs1_data_q\[5\] _01702_ _01703_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_72_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06573_ u_rf.reg6_q\[3\] _01555_ _01649_ u_rf.reg4_q\[3\] VGND VGND VPWR VPWR _01837_
+ sky130_fd_sc_hd__a22o_1
X_09361_ u_rf.reg2_q\[3\] _04434_ _04428_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08312_ u_rf.reg30_q\[7\] _03341_ _03342_ u_rf.reg10_q\[7\] _03508_ VGND VGND VPWR
+ VPWR _03509_ sky130_fd_sc_hd__a221o_1
X_09292_ _04385_ u_decod.rs2_data_q\[9\] _04386_ VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__and3_1
XANTENNA_12 _01605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _01763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08243_ _03436_ _03438_ _03440_ _03442_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_34 _03273_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 _03296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_56 _03353_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _03669_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _05271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _04827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08174_ _03364_ _03368_ _03372_ _03376_ VGND VGND VPWR VPWR _03377_ sky130_fd_sc_hd__or4_1
X_07125_ _01659_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__buf_6
XFILLER_0_140_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_50 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07056_ _01819_ _02300_ _01296_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__a21oi_1
Xoutput141 net141 VGND VGND VPWR VPWR icache_adr_o[16] sky130_fd_sc_hd__buf_4
Xoutput152 net152 VGND VGND VPWR VPWR icache_adr_o[26] sky130_fd_sc_hd__buf_4
XFILLER_0_113_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06007_ u_decod.rs2_data_q\[24\] u_decod.rs1_data_q\[24\] VGND VGND VPWR VPWR _01278_
+ sky130_fd_sc_hd__nand2_2
Xoutput130 net130 VGND VGND VPWR VPWR adr_o[7] sky130_fd_sc_hd__buf_2
Xoutput185 net185 VGND VGND VPWR VPWR store_data_o[26] sky130_fd_sc_hd__clkbuf_4
Xoutput163 net163 VGND VGND VPWR VPWR icache_adr_o[7] sky130_fd_sc_hd__clkbuf_4
Xoutput174 net174 VGND VGND VPWR VPWR store_data_o[16] sky130_fd_sc_hd__clkbuf_4
Xoutput196 net196 VGND VGND VPWR VPWR store_data_o[7] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_145_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07958_ _03164_ _03165_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[31\] sky130_fd_sc_hd__xor2_1
X_07889_ _02723_ _03048_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__nor2_1
X_06909_ u_rf.reg11_q\[10\] _01582_ _01665_ u_rf.reg8_q\[10\] VGND VGND VPWR VPWR
+ _02159_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09628_ u_rf.reg3_q\[18\] _04465_ _04582_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _04553_ VGND VGND VPWR VPWR _00082_ sky130_fd_sc_hd__clkbuf_1
X_12570_ clknet_leaf_64_clk _00607_ net346 VGND VGND VPWR VPWR u_rf.reg18_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11521_ _04738_ u_rf.reg30_q\[8\] _05621_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11452_ _05593_ VGND VGND VPWR VPWR _00935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10403_ _05036_ VGND VGND VPWR VPWR _00443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11383_ u_rf.reg28_q\[7\] net509 _05549_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__mux2_1
X_10334_ _04998_ VGND VGND VPWR VPWR _00412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ u_rf.reg12_q\[6\] _04951_ _04939_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__mux2_1
X_12004_ clknet_leaf_83_clk u_exe.bu_pc_res\[17\] net365 VGND VGND VPWR VPWR u_exe.pc_data_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10196_ _04899_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__buf_8
XFILLER_0_108_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_30_clk _00943_ net259 VGND VGND VPWR VPWR u_rf.reg29_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ clknet_leaf_123_clk _00874_ net231 VGND VGND VPWR VPWR u_rf.reg27_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12768_ clknet_leaf_119_clk _00805_ net249 VGND VGND VPWR VPWR u_rf.reg25_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12699_ clknet_leaf_12_clk _00736_ net243 VGND VGND VPWR VPWR u_rf.reg23_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_11719_ clknet_leaf_140_clk _00011_ net202 VGND VGND VPWR VPWR u_rf.reg2_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput21 icache_instr_i[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_1
Xinput10 icache_instr_i[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
XFILLER_0_37_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput32 icache_instr_i[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 load_data_i[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput54 load_data_i[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput76 reset_adr_i[1] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
Xinput65 reset_adr_i[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
Xinput87 reset_adr_i[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XFILLER_0_4_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_666 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08930_ _04074_ _04077_ _04081_ _04088_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08861_ _03998_ _04029_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__nor2_1
X_07812_ u_rf.reg12_q\[28\] _01610_ _02368_ u_rf.reg26_q\[28\] _03025_ VGND VGND VPWR
+ VPWR _03026_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_127_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08792_ u_rf.reg9_q\[29\] _03212_ _03295_ u_rf.reg20_q\[29\] VGND VGND VPWR VPWR
+ _03967_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07743_ _01472_ _02785_ _01500_ VGND VGND VPWR VPWR _02960_ sky130_fd_sc_hd__o21ai_1
X_07674_ u_rf.reg22_q\[25\] _01652_ _01673_ u_rf.reg2_q\[25\] VGND VGND VPWR VPWR
+ _02894_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_140_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09413_ _04427_ VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06625_ u_rf.reg11_q\[4\] _01583_ _01666_ u_rf.reg8_q\[4\] _01886_ VGND VGND VPWR
+ VPWR _01887_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09344_ u_decod.rf_ff_res_data_i\[0\] VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__buf_2
X_06556_ _01320_ _01763_ _01820_ _01312_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09275_ _01481_ _03998_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__nor2_1
XFILLER_0_75_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06487_ u_decod.rs1_data_q\[17\] _01446_ _01753_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_43_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08226_ u_rf.reg15_q\[3\] _03301_ _03303_ u_rf.reg24_q\[3\] _03426_ VGND VGND VPWR
+ VPWR _03427_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_758 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08157_ u_rf.reg22_q\[1\] _03275_ _03277_ u_rf.reg3_q\[1\] VGND VGND VPWR VPWR _03360_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07108_ _02345_ _02350_ _01757_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08088_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_655 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07039_ u_decod.pc_q_o\[12\] u_decod.pc_q_o\[13\] _02185_ VGND VGND VPWR VPWR _02284_
+ sky130_fd_sc_hd__and3_2
X_10050_ _04833_ VGND VGND VPWR VPWR _00293_ sky130_fd_sc_hd__clkbuf_1
X_10952_ _05328_ VGND VGND VPWR VPWR _00700_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10883_ _05291_ VGND VGND VPWR VPWR _00668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12622_ clknet_leaf_28_clk _00659_ net258 VGND VGND VPWR VPWR u_rf.reg20_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12553_ clknet_leaf_22_clk _00590_ net284 VGND VGND VPWR VPWR u_rf.reg18_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11504_ _05620_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__buf_6
XFILLER_0_108_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ clknet_leaf_111_clk _00521_ net316 VGND VGND VPWR VPWR u_rf.reg16_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11435_ _01534_ _04424_ _04936_ _05113_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__or4_4
XFILLER_0_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_780 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11366_ _05547_ VGND VGND VPWR VPWR _00895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10317_ u_decod.rf_ff_res_data_i\[23\] VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__buf_2
X_11297_ u_rf.reg26_q\[31\] u_decod.rf_ff_res_data_i\[31\] _05476_ VGND VGND VPWR
+ VPWR _05511_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10248_ _04940_ VGND VGND VPWR VPWR _00384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ _04902_ VGND VGND VPWR VPWR _00353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06410_ _01679_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07390_ _01057_ VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06341_ _01572_ _01551_ _01558_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__and3_4
XFILLER_0_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09060_ _04197_ _04198_ _04199_ _04200_ _04201_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[0\]
+ sky130_fd_sc_hd__a32o_1
X_06272_ u_decod.rf_ff_rd_adr_q_i\[1\] VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08011_ _03188_ _03198_ _03204_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__and3_4
XFILLER_0_123_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09962_ _04784_ u_rf.reg7_q\[30\] _04721_ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_430 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08913_ _04072_ _04073_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09893_ u_decod.rf_ff_res_data_i\[8\] VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08844_ u_decod.rs1_data_q\[3\] u_decod.branch_imm_q_o\[3\] VGND VGND VPWR VPWR _04015_
+ sky130_fd_sc_hd__and2_1
X_08775_ u_rf.reg28_q\[28\] _03556_ _03557_ u_rf.reg2_q\[28\] VGND VGND VPWR VPWR
+ _03951_ sky130_fd_sc_hd__a22o_1
X_05987_ u_decod.instr_unit_q\[0\] _01056_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__and2_1
X_07726_ u_rf.reg0_q\[26\] _01663_ _01674_ u_rf.reg2_q\[26\] VGND VGND VPWR VPWR _02944_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_255 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ _01430_ _01275_ _01277_ u_decod.instr_operation_q\[3\] _02877_ VGND VGND
+ VPWR VPWR _02878_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07588_ u_decod.rf_ff_res_data_i\[23\] _02358_ _02743_ _02792_ _02811_ VGND VGND
+ VPWR VPWR _02812_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06608_ _01808_ _01870_ _01423_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09327_ _04412_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_1
XFILLER_0_91_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06539_ net201 _01804_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_153_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09258_ _04160_ _04206_ _04197_ _04371_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[28\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09189_ u_decod.pc_q_o\[19\] u_decod.branch_imm_q_o\[19\] VGND VGND VPWR VPWR _04312_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08209_ _03219_ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__buf_8
XFILLER_0_43_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11220_ _05470_ VGND VGND VPWR VPWR _00826_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11151_ u_rf.reg24_q\[26\] _04993_ _05427_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__mux2_1
X_10102_ _04860_ VGND VGND VPWR VPWR _00318_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11082_ _05397_ VGND VGND VPWR VPWR _00761_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10033_ _04823_ VGND VGND VPWR VPWR _00286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11984_ clknet_leaf_103_clk u_decod.dec0.is_shift net335 VGND VGND VPWR VPWR u_decod.instr_unit_q\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_10935_ u_rf.reg21_q\[20\] _04980_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10866_ u_rf.reg20_q\[20\] _04980_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12605_ clknet_leaf_15_clk _00642_ net246 VGND VGND VPWR VPWR u_rf.reg20_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10797_ _05223_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__buf_6
XFILLER_0_38_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12536_ clknet_leaf_67_clk _00573_ net349 VGND VGND VPWR VPWR u_rf.reg17_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12467_ clknet_leaf_52_clk _00504_ net305 VGND VGND VPWR VPWR u_rf.reg15_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11418_ _05575_ VGND VGND VPWR VPWR _00919_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_840 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12398_ clknet_leaf_27_clk _00435_ net258 VGND VGND VPWR VPWR u_rf.reg13_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11349_ _04770_ u_rf.reg27_q\[23\] _05535_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_783 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06890_ _01302_ _01702_ _01703_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__o21a_1
X_05910_ u_decod.dec0.instr_i\[1\] u_decod.dec0.instr_i\[3\] u_decod.dec0.instr_i\[2\]
+ _01198_ _01199_ VGND VGND VPWR VPWR _01200_ sky130_fd_sc_hd__a41o_1
X_05841_ u_decod.pc0_q_i\[15\] _01143_ VGND VGND VPWR VPWR _01148_ sky130_fd_sc_hd__nand2_1
X_08560_ u_rf.reg25_q\[18\] _03315_ _03325_ u_rf.reg5_q\[18\] _03745_ VGND VGND VPWR
+ VPWR _03746_ sky130_fd_sc_hd__a221o_1
X_05772_ _01074_ _01092_ _01094_ VGND VGND VPWR VPWR _01095_ sky130_fd_sc_hd__and3_1
X_07511_ _01359_ _01395_ _02674_ _01374_ _01396_ VGND VGND VPWR VPWR _02738_ sky130_fd_sc_hd__a311o_1
X_08491_ u_rf.reg1_q\[15\] _03310_ _03312_ u_rf.reg14_q\[15\] VGND VGND VPWR VPWR
+ _03680_ sky130_fd_sc_hd__a22o_1
X_07442_ _02572_ _02573_ _02616_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__and3_1
X_07373_ u_rf.reg0_q\[19\] _01662_ _01597_ u_rf.reg13_q\[19\] VGND VGND VPWR VPWR
+ _02605_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09112_ _04244_ _04245_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06324_ _01593_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_40_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06255_ _01520_ u_decod.exe_ff_rd_adr_q_i\[0\] u_decod.exe_ff_rd_adr_q_i\[2\] _01522_
+ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09043_ _01325_ _01326_ _01311_ _01316_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_588 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06186_ _01450_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09945_ _04773_ VGND VGND VPWR VPWR _00248_ sky130_fd_sc_hd__clkbuf_1
X_09876_ _04726_ u_rf.reg7_q\[2\] _04722_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ u_decod.branch_imm_q_o\[0\] _01061_ _01060_ _03999_ VGND VGND VPWR VPWR _04000_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ u_decod.exe_ff_res_data_i\[27\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[27\]
+ _03934_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__a221o_1
X_08689_ u_rf.reg6_q\[24\] _03387_ _03388_ u_rf.reg13_q\[24\] VGND VGND VPWR VPWR
+ _03869_ sky130_fd_sc_hd__a22o_1
X_07709_ _01260_ _02916_ _02927_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_726 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10720_ _05205_ VGND VGND VPWR VPWR _00591_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10651_ u_rf.reg17_q\[15\] _04970_ _05163_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10582_ _05132_ VGND VGND VPWR VPWR _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12321_ clknet_leaf_118_clk _00358_ net326 VGND VGND VPWR VPWR u_rf.reg11_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12252_ clknet_leaf_128_clk _00289_ net234 VGND VGND VPWR VPWR u_rf.reg9_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11203_ _05461_ VGND VGND VPWR VPWR _00818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12183_ clknet_leaf_50_clk _00220_ net352 VGND VGND VPWR VPWR u_rf.reg6_q\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_71_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ u_rf.reg24_q\[18\] _04976_ _05416_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__mux2_1
X_11065_ _05388_ VGND VGND VPWR VPWR _00753_ sky130_fd_sc_hd__clkbuf_1
X_10016_ u_rf.reg8_q\[22\] _04474_ _04812_ VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11967_ clknet_leaf_83_clk net453 net365 VGND VGND VPWR VPWR u_decod.pc_q_o\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_102_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_86_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10918_ u_rf.reg21_q\[12\] _04964_ _05308_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_444 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11898_ clknet_leaf_96_clk u_decod.rs2_data_nxt\[19\] net333 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10849_ u_rf.reg20_q\[12\] _04964_ _05271_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12519_ clknet_leaf_4_clk _00556_ net212 VGND VGND VPWR VPWR u_rf.reg17_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06040_ _01309_ _01310_ VGND VGND VPWR VPWR _01311_ sky130_fd_sc_hd__or2b_2
XFILLER_0_140_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07991_ _03187_ _03196_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__nor2_2
Xfanout219 net220 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
Xfanout208 net210 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ _04646_ VGND VGND VPWR VPWR _04647_ sky130_fd_sc_hd__buf_6
X_06942_ u_decod.rs1_data_q\[26\] _01454_ _01753_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09661_ _04609_ VGND VGND VPWR VPWR _00128_ sky130_fd_sc_hd__clkbuf_1
X_06873_ u_rf.reg6_q\[9\] _01554_ _01651_ u_rf.reg22_q\[9\] VGND VGND VPWR VPWR _02125_
+ sky130_fd_sc_hd__a22o_1
X_08612_ u_rf.reg22_q\[21\] _03274_ _03410_ u_rf.reg3_q\[21\] VGND VGND VPWR VPWR
+ _03795_ sky130_fd_sc_hd__a22o_1
X_05824_ _01133_ _01106_ _01134_ VGND VGND VPWR VPWR _01135_ sky130_fd_sc_hd__and3b_1
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09592_ _04572_ VGND VGND VPWR VPWR _00096_ sky130_fd_sc_hd__clkbuf_1
X_08543_ u_decod.rf_ff_res_data_i\[17\] _03382_ _03729_ _03404_ VGND VGND VPWR VPWR
+ _03730_ sky130_fd_sc_hd__a22o_1
X_05755_ _01076_ _01077_ VGND VGND VPWR VPWR _01078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08474_ u_rf.reg7_q\[14\] _03314_ _03315_ u_rf.reg25_q\[14\] _03663_ VGND VGND VPWR
+ VPWR _03664_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_137_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ u_rf.reg30_q\[20\] _01580_ _01625_ u_rf.reg28_q\[20\] VGND VGND VPWR VPWR
+ _02655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07356_ _01377_ _01431_ _01434_ _02588_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07287_ u_rf.reg30_q\[17\] _01579_ _01591_ u_rf.reg18_q\[17\] VGND VGND VPWR VPWR
+ _02523_ sky130_fd_sc_hd__a22o_1
X_06307_ _01522_ _01537_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_188 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09026_ net133 _04170_ VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06238_ u_decod.pc_q_o\[0\] _01485_ _01492_ _01059_ _01508_ VGND VGND VPWR VPWR _01509_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06169_ u_decod.instr_operation_q\[4\] _01420_ _01421_ _01426_ _01439_ VGND VGND
+ VPWR VPWR _01440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09928_ _04761_ u_rf.reg7_q\[19\] _04743_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09859_ _04715_ VGND VGND VPWR VPWR _00220_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ clknet_leaf_3_clk _00907_ net213 VGND VGND VPWR VPWR u_rf.reg28_q\[11\] sky130_fd_sc_hd__dfrtp_1
X_11821_ clknet_leaf_94_clk net8 net339 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_102 _05632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net469 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 u_decod.rs1_data_q\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _01679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _04874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_168 u_decod.pc_q_o\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11752_ clknet_leaf_3_clk _00044_ net211 VGND VGND VPWR VPWR u_rf.reg1_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11683_ u_decod.branch_imm_q_o\[20\] _02647_ _05696_ VGND VGND VPWR VPWR _05716_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _05196_ VGND VGND VPWR VPWR _00583_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_81_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10634_ u_rf.reg17_q\[7\] _04953_ _05152_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_864 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12304_ clknet_leaf_34_clk _00341_ net268 VGND VGND VPWR VPWR u_rf.reg10_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ _05123_ VGND VGND VPWR VPWR _00518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10496_ _04736_ u_rf.reg15_q\[7\] _05078_ VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__mux2_1
X_12235_ clknet_leaf_1_clk _00272_ net221 VGND VGND VPWR VPWR u_rf.reg8_q\[16\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12166_ clknet_leaf_139_clk _00203_ net202 VGND VGND VPWR VPWR u_rf.reg6_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ _05404_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__buf_8
X_12097_ clknet_leaf_119_clk _00134_ net250 VGND VGND VPWR VPWR u_rf.reg4_q\[6\] sky130_fd_sc_hd__dfrtp_1
Xinput8 icache_instr_i[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
X_11048_ _05379_ VGND VGND VPWR VPWR _00745_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12999_ clknet_leaf_91_clk _01036_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[12\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_157_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08190_ u_rf.reg27_q\[2\] _03318_ _03320_ u_rf.reg19_q\[2\] _03391_ VGND VGND VPWR
+ VPWR _03392_ sky130_fd_sc_hd__a221o_1
X_07210_ _01388_ u_decod.rs1_data_q\[8\] _01061_ _01747_ _01455_ _01461_ VGND VGND
+ VPWR VPWR _02449_ sky130_fd_sc_hd__mux4_2
XFILLER_0_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07141_ u_rf.reg1_q\[14\] _01587_ _01667_ u_rf.reg8_q\[14\] VGND VGND VPWR VPWR _02383_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07072_ u_rf.reg5_q\[13\] _01568_ _01555_ u_rf.reg6_q\[13\] VGND VGND VPWR VPWR _02316_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06023_ _01291_ _01293_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07974_ u_decod.dec0.instr_i\[15\] VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__inv_2
X_09713_ _04636_ VGND VGND VPWR VPWR _00153_ sky130_fd_sc_hd__clkbuf_1
X_06925_ _02165_ _02174_ _01678_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__o21a_1
X_09644_ _04599_ VGND VGND VPWR VPWR _00121_ sky130_fd_sc_hd__clkbuf_1
X_06856_ u_decod.pc_q_o\[9\] _02054_ _02108_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__o21ai_1
X_05807_ u_decod.pc0_q_i\[6\] net382 u_decod.pc0_q_i\[7\] VGND VGND VPWR VPWR _01122_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_143_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ u_rf.reg0_q\[26\] _04482_ _04555_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06787_ u_decod.rs1_data_q\[8\] _01445_ _01494_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08526_ u_rf.reg31_q\[17\] _03210_ _03211_ u_rf.reg11_q\[17\] VGND VGND VPWR VPWR
+ _03713_ sky130_fd_sc_hd__a22o_1
X_05738_ _01058_ _01063_ VGND VGND VPWR VPWR _01064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_37_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_718 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08457_ net450 _03565_ _03647_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07408_ u_decod.pc_q_o\[20\] _02578_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08388_ u_rf.reg0_q\[10\] _03176_ _03329_ u_rf.reg12_q\[10\] _03581_ VGND VGND VPWR
+ VPWR _03582_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_823 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07339_ _02486_ _02530_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10350_ _04726_ u_rf.reg13_q\[2\] _05006_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09009_ _04135_ _04152_ _04155_ VGND VGND VPWR VPWR _04156_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10281_ u_rf.reg12_q\[11\] _04962_ _04960_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__mux2_1
X_12020_ clknet_leaf_98_clk u_decod.exe_ff_res_data_i\[0\] net330 VGND VGND VPWR VPWR
+ u_decod.rf_ff_res_data_i\[0\] sky130_fd_sc_hd__dfrtp_4
X_12922_ clknet_leaf_94_clk _00959_ net339 VGND VGND VPWR VPWR u_rf.reg29_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
X_12853_ clknet_leaf_47_clk _00890_ net299 VGND VGND VPWR VPWR u_rf.reg27_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ clknet_leaf_36_clk _00821_ net271 VGND VGND VPWR VPWR u_rf.reg25_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11804_ clknet_leaf_81_clk net158 net361 VGND VGND VPWR VPWR u_decod.pc0_q_i\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11735_ clknet_leaf_51_clk _00027_ net307 VGND VGND VPWR VPWR u_rf.reg2_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_835 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11666_ _05707_ VGND VGND VPWR VPWR _01035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_378 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10617_ _05150_ VGND VGND VPWR VPWR _00543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11597_ _05670_ VGND VGND VPWR VPWR _01003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10548_ u_decod.rf_ff_rd_adr_q_i\[4\] u_decod.rf_write_v_q_i VGND VGND VPWR VPWR
+ _05113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10479_ _05076_ VGND VGND VPWR VPWR _00479_ sky130_fd_sc_hd__clkbuf_1
X_12218_ clknet_leaf_94_clk _00255_ net339 VGND VGND VPWR VPWR u_rf.reg7_q\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12149_ clknet_leaf_46_clk _00186_ net298 VGND VGND VPWR VPWR u_rf.reg5_q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06710_ _01968_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[6\] sky130_fd_sc_hd__inv_2
X_07690_ u_decod.pc_q_o\[26\] _02868_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__and2_1
X_06641_ _01311_ _01323_ _01860_ _01765_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06572_ u_rf.reg3_q\[3\] _01605_ _01631_ u_rf.reg17_q\[3\] _01835_ VGND VGND VPWR
+ VPWR _01836_ sky130_fd_sc_hd__a221o_1
X_09360_ u_decod.rf_ff_res_data_i\[3\] VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__buf_2
XFILLER_0_157_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08311_ u_rf.reg26_q\[7\] _03344_ _03345_ u_rf.reg21_q\[7\] VGND VGND VPWR VPWR _03508_
+ sky130_fd_sc_hd__a22o_1
X_09291_ _04392_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_1
XFILLER_0_129_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_13 _01615_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08242_ u_rf.reg31_q\[4\] _03290_ _03292_ u_rf.reg11_q\[4\] _03441_ VGND VGND VPWR
+ VPWR _03442_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _03305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_57 _03356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _01772_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_68 _03670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_79 _04838_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08173_ u_rf.reg15_q\[1\] _03373_ _03374_ u_rf.reg24_q\[1\] _03375_ VGND VGND VPWR
+ VPWR _03376_ sky130_fd_sc_hd__a221o_1
X_07124_ u_rf.reg3_q\[14\] _02363_ _02364_ u_rf.reg21_q\[14\] _02365_ VGND VGND VPWR
+ VPWR _02366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_62 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07055_ _01295_ _01697_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput120 net120 VGND VGND VPWR VPWR adr_o[27] sky130_fd_sc_hd__clkbuf_4
Xoutput142 net142 VGND VGND VPWR VPWR icache_adr_o[17] sky130_fd_sc_hd__buf_2
XFILLER_0_140_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06006_ _01275_ _01276_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__and2_2
XFILLER_0_101_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput131 net131 VGND VGND VPWR VPWR adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput153 net153 VGND VGND VPWR VPWR icache_adr_o[27] sky130_fd_sc_hd__clkbuf_4
Xoutput186 net186 VGND VGND VPWR VPWR store_data_o[27] sky130_fd_sc_hd__clkbuf_4
Xoutput164 net164 VGND VGND VPWR VPWR icache_adr_o[8] sky130_fd_sc_hd__buf_4
Xoutput175 net175 VGND VGND VPWR VPWR store_data_o[17] sky130_fd_sc_hd__clkbuf_4
Xoutput197 net197 VGND VGND VPWR VPWR store_data_o[8] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07957_ _03041_ _03042_ _03081_ _03126_ _01897_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__o41a_1
X_06908_ u_rf.reg23_q\[10\] _01611_ _01655_ u_rf.reg10_q\[10\] _02157_ VGND VGND VPWR
+ VPWR _02158_ sky130_fd_sc_hd__a221o_1
X_07888_ _01502_ _03009_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09627_ _04590_ VGND VGND VPWR VPWR _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06839_ _02091_ _01337_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09558_ u_rf.reg0_q\[18\] _04465_ _04544_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08509_ u_rf.reg9_q\[16\] _03294_ _03296_ u_rf.reg20_q\[16\] VGND VGND VPWR VPWR
+ _03697_ sky130_fd_sc_hd__a22o_1
X_09489_ u_rf.reg1_q\[18\] _04465_ _04507_ VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _05629_ VGND VGND VPWR VPWR _00967_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11451_ _04736_ u_rf.reg29_q\[7\] _05585_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10402_ _04778_ u_rf.reg13_q\[27\] _05028_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__mux2_1
X_11382_ _05556_ VGND VGND VPWR VPWR _00902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10333_ u_rf.reg12_q\[28\] _04997_ _04981_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ u_decod.rf_ff_res_data_i\[6\] VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__buf_2
X_12003_ clknet_leaf_83_clk u_exe.bu_pc_res\[16\] net366 VGND VGND VPWR VPWR u_exe.pc_data_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10195_ _04910_ VGND VGND VPWR VPWR _00361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ clknet_leaf_24_clk _00942_ net267 VGND VGND VPWR VPWR u_rf.reg29_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ clknet_leaf_111_clk _00873_ net316 VGND VGND VPWR VPWR u_rf.reg27_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12767_ clknet_leaf_132_clk _00804_ net228 VGND VGND VPWR VPWR u_rf.reg25_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12698_ clknet_leaf_94_clk _00735_ net339 VGND VGND VPWR VPWR u_rf.reg22_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11718_ clknet_leaf_121_clk _00010_ net247 VGND VGND VPWR VPWR u_rf.reg2_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11649_ _05698_ VGND VGND VPWR VPWR _01027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 icache_instr_i[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 icache_instr_i[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
XFILLER_0_142_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_480 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput55 load_data_i[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_1
Xinput44 load_data_i[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput33 load_data_i[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput77 reset_adr_i[20] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
Xinput88 reset_adr_i[30] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
Xinput66 reset_adr_i[10] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08860_ _04025_ net380 VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__xnor2_1
X_07811_ u_rf.reg19_q\[28\] _02665_ _02697_ u_rf.reg4_q\[28\] VGND VGND VPWR VPWR
+ _03025_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08791_ u_rf.reg15_q\[29\] _03300_ _03328_ u_rf.reg12_q\[29\] _03965_ VGND VGND VPWR
+ VPWR _03966_ sky130_fd_sc_hd__a221o_1
X_07742_ _02619_ net52 _02618_ VGND VGND VPWR VPWR _02959_ sky130_fd_sc_hd__a21bo_1
X_07673_ _02886_ _02888_ _02890_ _02892_ VGND VGND VPWR VPWR _02893_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_140_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ u_decod.rf_ff_res_data_i\[20\] VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06624_ u_rf.reg1_q\[4\] _01586_ _01635_ u_rf.reg9_q\[4\] VGND VGND VPWR VPWR _01886_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09343_ _04420_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_1
XFILLER_0_59_150 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06555_ _01819_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__buf_4
X_09274_ _04197_ _04383_ _04384_ _04200_ _04174_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[31\]
+ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_43_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06486_ _01494_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08225_ u_rf.reg6_q\[3\] _03387_ _03388_ u_rf.reg13_q\[3\] VGND VGND VPWR VPWR _03426_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08156_ u_rf.reg18_q\[1\] _03353_ _03355_ u_rf.reg23_q\[1\] _03358_ VGND VGND VPWR
+ VPWR _03359_ sky130_fd_sc_hd__a221o_1
X_07107_ _01464_ _02347_ _02349_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__a21oi_1
X_08087_ _03211_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07038_ _02281_ _01347_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08989_ _04137_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10951_ u_rf.reg21_q\[28\] _04997_ _05319_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10882_ u_rf.reg20_q\[28\] _04997_ _05282_ VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12621_ clknet_leaf_5_clk _00658_ net217 VGND VGND VPWR VPWR u_rf.reg20_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12552_ clknet_leaf_18_clk _00589_ net288 VGND VGND VPWR VPWR u_rf.reg18_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_304 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11503_ _04425_ _04936_ _05114_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__or3_4
XFILLER_0_65_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12483_ clknet_leaf_109_clk _00520_ net313 VGND VGND VPWR VPWR u_rf.reg16_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11434_ _05583_ VGND VGND VPWR VPWR _00927_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_91_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_792 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11365_ _04786_ u_rf.reg27_q\[31\] _05512_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_100_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_100_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_245 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10316_ _04986_ VGND VGND VPWR VPWR _00406_ sky130_fd_sc_hd__clkbuf_1
X_11296_ _05510_ VGND VGND VPWR VPWR _00862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10247_ u_rf.reg12_q\[0\] _04935_ _04939_ VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ _04724_ u_rf.reg11_q\[1\] _04900_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12819_ clknet_leaf_66_clk _00856_ net356 VGND VGND VPWR VPWR u_rf.reg26_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_542 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06340_ _01609_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__buf_6
X_06271_ _01534_ u_decod.dec0.instr_i\[20\] u_decod.dec0.instr_i\[23\] _01535_ _01540_
+ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_586 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08010_ _03171_ _03172_ _03201_ VGND VGND VPWR VPWR _03216_ sky130_fd_sc_hd__and3_2
XFILLER_0_72_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_442 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09961_ u_decod.rf_ff_res_data_i\[30\] VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__buf_2
XFILLER_0_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08912_ _01292_ u_decod.branch_imm_q_o\[14\] VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_139_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09892_ _04737_ VGND VGND VPWR VPWR _00231_ sky130_fd_sc_hd__clkbuf_1
X_08843_ _04012_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__and2_1
X_08774_ u_rf.reg27_q\[28\] _03365_ _03366_ u_rf.reg19_q\[28\] _03949_ VGND VGND VPWR
+ VPWR _03950_ sky130_fd_sc_hd__a221o_1
X_05986_ net463 VGND VGND VPWR VPWR u_decod.exe_ff_write_v_q_i sky130_fd_sc_hd__inv_2
XFILLER_0_33_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07725_ u_rf.reg22_q\[26\] _01654_ _01668_ u_rf.reg8_q\[26\] _02942_ VGND VGND VPWR
+ VPWR _02943_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07656_ u_decod.rs2_data_q\[25\] u_decod.rs1_data_q\[25\] _02781_ VGND VGND VPWR
+ VPWR _02877_ sky130_fd_sc_hd__and3_1
X_07587_ _02794_ _02801_ _02810_ _02359_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__o31a_2
XFILLER_0_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06607_ _01756_ _01869_ _01688_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09326_ _04409_ u_decod.rs2_data_q\[24\] _04410_ VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06538_ _01511_ _01528_ _01682_ _01803_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09257_ _04367_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08208_ _03218_ VGND VGND VPWR VPWR _03409_ sky130_fd_sc_hd__buf_6
X_06469_ _01713_ u_decod.exe_ff_res_data_i\[1\] _01717_ _01736_ VGND VGND VPWR VPWR
+ _01737_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_153_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09188_ u_decod.pc_q_o\[19\] u_decod.branch_imm_q_o\[19\] VGND VGND VPWR VPWR _04311_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08139_ _03282_ VGND VGND VPWR VPWR _03342_ sky130_fd_sc_hd__buf_6
X_11150_ _05433_ VGND VGND VPWR VPWR _00793_ sky130_fd_sc_hd__clkbuf_1
X_10101_ u_rf.reg9_q\[30\] _04490_ _04826_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11081_ _04774_ u_rf.reg23_q\[25\] _05391_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ u_rf.reg8_q\[30\] _04490_ _04789_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__mux2_1
X_11983_ clknet_leaf_103_clk u_decod.dec0.is_arithm net335 VGND VGND VPWR VPWR u_decod.instr_unit_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10934_ _05296_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_104_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10865_ _05259_ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_27_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12604_ clknet_leaf_127_clk _00641_ net235 VGND VGND VPWR VPWR u_rf.reg20_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12535_ clknet_leaf_71_clk _00572_ net353 VGND VGND VPWR VPWR u_rf.reg17_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10796_ _05245_ VGND VGND VPWR VPWR _00627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12466_ clknet_leaf_39_clk _00503_ net277 VGND VGND VPWR VPWR u_rf.reg15_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11417_ u_rf.reg28_q\[23\] u_decod.rf_ff_res_data_i\[23\] _05571_ VGND VGND VPWR
+ VPWR _05575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12397_ clknet_leaf_7_clk _00434_ net217 VGND VGND VPWR VPWR u_rf.reg13_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11348_ _05538_ VGND VGND VPWR VPWR _00886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11279_ u_rf.reg26_q\[22\] u_decod.rf_ff_res_data_i\[22\] _05499_ VGND VGND VPWR
+ VPWR _05502_ sky130_fd_sc_hd__mux2_1
X_13018_ clknet_leaf_65_clk _01055_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[31\]
+ sky130_fd_sc_hd__dfxtp_1
X_05840_ u_decod.pc0_q_i\[15\] _01143_ VGND VGND VPWR VPWR _01147_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07510_ _01372_ _01373_ _01361_ _02637_ _01397_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__a221o_1
X_05771_ _01076_ _01093_ VGND VGND VPWR VPWR _01094_ sky130_fd_sc_hd__and2_1
X_08490_ _03672_ _03674_ _03676_ _03678_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__or4_1
XFILLER_0_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_418 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07441_ _02357_ u_decod.exe_ff_res_data_i\[20\] _02670_ VGND VGND VPWR VPWR _02671_
+ sky130_fd_sc_hd__a21o_1
X_07372_ _01586_ VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__buf_6
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09111_ u_decod.pc_q_o\[8\] u_decod.branch_imm_q_o\[8\] VGND VGND VPWR VPWR _04245_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06323_ _01572_ _01515_ _01558_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__and3_2
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09042_ _01263_ _01270_ _04183_ _04184_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__or4_4
X_06254_ _01520_ u_decod.exe_ff_rd_adr_q_i\[0\] u_decod.exe_ff_rd_adr_q_i\[4\] _01512_
+ _01523_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06185_ net376 _01380_ u_decod.rs1_data_q\[9\] u_decod.rs1_data_q\[25\] _01454_ _01455_
+ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_147_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09944_ _04772_ u_rf.reg7_q\[24\] _04764_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09875_ u_decod.rf_ff_res_data_i\[2\] VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_5_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ u_decod.branch_imm_q_o\[1\] net375 VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _03924_ _03933_ _03378_ VGND VGND VPWR VPWR _03934_ sky130_fd_sc_hd__o21a_1
X_05969_ u_decod.dec0.instr_i\[5\] _01076_ _01086_ _01093_ VGND VGND VPWR VPWR _01246_
+ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_156_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08688_ u_rf.reg27_q\[24\] _03365_ _03366_ u_rf.reg19_q\[24\] _03867_ VGND VGND VPWR
+ VPWR _03868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07708_ _01746_ _02920_ _02924_ _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07639_ u_decod.rf_ff_res_data_i\[24\] _02358_ _02743_ _02841_ _02860_ VGND VGND
+ VPWR VPWR _02861_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_95_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10650_ _05168_ VGND VGND VPWR VPWR _00558_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09309_ _04402_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_146_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10581_ u_rf.reg16_q\[14\] _04968_ _05127_ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12320_ clknet_leaf_117_clk _00357_ net323 VGND VGND VPWR VPWR u_rf.reg11_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12251_ clknet_leaf_122_clk _00288_ net241 VGND VGND VPWR VPWR u_rf.reg9_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11202_ u_rf.reg25_q\[18\] _04976_ _05452_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_1
X_12182_ clknet_leaf_48_clk _00219_ net306 VGND VGND VPWR VPWR u_rf.reg6_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_250 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11133_ _05424_ VGND VGND VPWR VPWR _00785_ sky130_fd_sc_hd__clkbuf_1
X_11064_ _04757_ u_rf.reg23_q\[17\] _05380_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__mux2_1
X_10015_ _04814_ VGND VGND VPWR VPWR _00277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11966_ clknet_leaf_82_clk net462 net361 VGND VGND VPWR VPWR u_decod.pc_q_o\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_86_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10917_ _05310_ VGND VGND VPWR VPWR _00683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11897_ clknet_leaf_96_clk u_decod.rs2_data_nxt\[18\] net333 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10848_ _05273_ VGND VGND VPWR VPWR _00651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10779_ u_rf.reg19_q\[11\] _04962_ _05235_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12518_ clknet_leaf_139_clk _00555_ net203 VGND VGND VPWR VPWR u_rf.reg17_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12449_ clknet_leaf_117_clk _00486_ net326 VGND VGND VPWR VPWR u_rf.reg15_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_256 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07990_ _01539_ _03188_ _03189_ _03195_ VGND VGND VPWR VPWR _03196_ sky130_fd_sc_hd__a211o_1
Xfanout209 net210 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_4
X_06941_ u_decod.rs1_data_q\[18\] _01454_ _01753_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09660_ u_rf.reg4_q\[0\] _04421_ _04608_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__mux2_1
X_08611_ net445 _03773_ _03793_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[20\]
+ sky130_fd_sc_hd__a22o_1
X_06872_ u_rf.reg0_q\[9\] _01516_ _01599_ u_rf.reg15_q\[9\] _02123_ VGND VGND VPWR
+ VPWR _02124_ sky130_fd_sc_hd__a221o_1
X_05823_ u_decod.pc0_q_i\[11\] net394 VGND VGND VPWR VPWR _01134_ sky130_fd_sc_hd__or2_1
X_09591_ u_rf.reg3_q\[0\] _04421_ _04571_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__mux2_1
X_08542_ _03712_ _03719_ _03728_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__or3_2
X_05754_ u_decod.dec0.funct3\[2\] u_decod.dec0.instr_i\[0\] VGND VGND VPWR VPWR _01077_
+ sky130_fd_sc_hd__nand2b_1
X_08473_ u_rf.reg1_q\[14\] _03231_ _03232_ u_rf.reg14_q\[14\] VGND VGND VPWR VPWR
+ _03663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07424_ u_rf.reg23_q\[20\] _02652_ _01654_ u_rf.reg22_q\[20\] _02653_ VGND VGND VPWR
+ VPWR _02654_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07355_ _01377_ _01378_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07286_ u_rf.reg20_q\[17\] _01644_ _01670_ u_rf.reg27_q\[17\] _02521_ VGND VGND VPWR
+ VPWR _02522_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06306_ _01575_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_150_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09025_ _04168_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06237_ _01424_ _01503_ _01506_ _01507_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_595 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06168_ _01061_ _01425_ _01429_ _01432_ _01438_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__a311o_1
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06099_ _01368_ _01369_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09927_ u_decod.rf_ff_res_data_i\[19\] VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_148_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09858_ u_rf.reg6_q\[28\] _04486_ _04706_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__mux2_1
X_09789_ u_rf.reg5_q\[28\] _04486_ _04669_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__mux2_1
X_08809_ u_rf.reg22_q\[30\] _03274_ _03276_ u_rf.reg3_q\[30\] VGND VGND VPWR VPWR
+ _03983_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 _05668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11820_ clknet_leaf_93_clk net7 net339 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_125 net509 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 u_decod.rs1_data_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_147 _03310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_158 _05017_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _01716_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ clknet_leaf_4_clk _00043_ net202 VGND VGND VPWR VPWR u_rf.reg1_q\[11\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_80_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10702_ u_rf.reg18_q\[7\] _04953_ _05188_ VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__mux2_1
XANTENNA_169 u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_154_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11682_ _05715_ VGND VGND VPWR VPWR _01043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _05159_ VGND VGND VPWR VPWR _00550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10564_ u_rf.reg16_q\[6\] _04951_ _05116_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12303_ clknet_leaf_42_clk _00340_ net295 VGND VGND VPWR VPWR u_rf.reg10_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10495_ _05085_ VGND VGND VPWR VPWR _00486_ sky130_fd_sc_hd__clkbuf_1
X_12234_ clknet_leaf_29_clk _00271_ net257 VGND VGND VPWR VPWR u_rf.reg8_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12165_ clknet_leaf_122_clk _00202_ net241 VGND VGND VPWR VPWR u_rf.reg6_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_112_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11116_ _05415_ VGND VGND VPWR VPWR _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12096_ clknet_leaf_114_clk _00133_ net323 VGND VGND VPWR VPWR u_rf.reg4_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_11047_ _04740_ u_rf.reg23_q\[9\] _05369_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__mux2_1
Xinput9 icache_instr_i[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12998_ clknet_leaf_91_clk _01035_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[11\]
+ sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_71_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_412 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11949_ clknet_leaf_98_clk u_decod.dec0.rd_o\[3\] net331 VGND VGND VPWR VPWR u_decod.exe_ff_rd_adr_q_i\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07140_ u_rf.reg17_q\[14\] _02379_ _02380_ u_rf.reg10_q\[14\] _02381_ VGND VGND VPWR
+ VPWR _02382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07071_ u_rf.reg0_q\[13\] _01663_ _01636_ u_rf.reg9_q\[13\] _02314_ VGND VGND VPWR
+ VPWR _02315_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06022_ u_decod.rs2_data_q\[14\] _01292_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_387 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09712_ u_rf.reg4_q\[25\] _04480_ _04630_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__mux2_1
X_07973_ u_decod.dec0.instr_i\[18\] u_decod.exe_ff_rd_adr_q_i\[3\] VGND VGND VPWR
+ VPWR _03179_ sky130_fd_sc_hd__xor2_1
X_06924_ _02167_ _02169_ _02171_ _02173_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__or4_1
X_09643_ u_rf.reg3_q\[25\] _04480_ _04593_ VGND VGND VPWR VPWR _04599_ sky130_fd_sc_hd__mux2_1
X_06855_ u_decod.pc_q_o\[9\] _02054_ _01764_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__a21oi_1
X_09574_ _04561_ VGND VGND VPWR VPWR _00089_ sky130_fd_sc_hd__clkbuf_1
X_05806_ u_decod.pc0_q_i\[6\] u_decod.pc0_q_i\[7\] _01113_ VGND VGND VPWR VPWR _01121_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_143_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08525_ u_rf.reg30_q\[17\] _03341_ _03342_ u_rf.reg10_q\[17\] _03711_ VGND VGND VPWR
+ VPWR _03712_ sky130_fd_sc_hd__a221o_1
X_06786_ _01996_ _02040_ _01422_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_62_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
X_05737_ net393 _01062_ VGND VGND VPWR VPWR _01063_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08456_ u_decod.exe_ff_res_data_i\[13\] _03381_ _03646_ VGND VGND VPWR VPWR _03647_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_426 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07407_ u_decod.pc_q_o\[20\] _02578_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ u_rf.reg28_q\[10\] _03331_ _03333_ u_rf.reg2_q\[10\] VGND VGND VPWR VPWR
+ _03581_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07338_ _01772_ u_decod.exe_ff_res_data_i\[18\] _02571_ VGND VGND VPWR VPWR _02572_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07269_ u_decod.pc_q_o\[15\] u_decod.pc_q_o\[16\] u_decod.pc_q_o\[17\] _02335_ VGND
+ VGND VPWR VPWR _02506_ sky130_fd_sc_hd__and4_1
XFILLER_0_104_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09008_ _04138_ _04144_ _04153_ _04149_ _04154_ VGND VGND VPWR VPWR _04155_ sky130_fd_sc_hd__o41a_1
XFILLER_0_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10280_ u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__buf_2
XFILLER_0_131_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12921_ clknet_leaf_63_clk _00958_ net342 VGND VGND VPWR VPWR u_rf.reg29_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12852_ clknet_leaf_31_clk _00889_ net264 VGND VGND VPWR VPWR u_rf.reg27_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12783_ clknet_leaf_37_clk _00820_ net272 VGND VGND VPWR VPWR u_rf.reg25_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_53_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
X_11803_ clknet_leaf_81_clk net157 net368 VGND VGND VPWR VPWR u_decod.pc0_q_i\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11734_ clknet_leaf_44_clk _00026_ net296 VGND VGND VPWR VPWR u_rf.reg2_q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11665_ u_decod.branch_imm_q_o\[11\] _02204_ _05696_ VGND VGND VPWR VPWR _05707_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_10616_ u_rf.reg16_q\[31\] _05003_ _05115_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_733 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11596_ _04745_ u_rf.reg31_q\[11\] _05668_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10547_ _05112_ VGND VGND VPWR VPWR _00511_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10478_ _04786_ u_rf.reg14_q\[31\] _05041_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12217_ clknet_leaf_57_clk _00254_ net292 VGND VGND VPWR VPWR u_rf.reg7_q\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12148_ clknet_leaf_32_clk _00185_ net262 VGND VGND VPWR VPWR u_rf.reg5_q\[25\] sky130_fd_sc_hd__dfrtp_1
X_12079_ clknet_leaf_35_clk _00116_ net272 VGND VGND VPWR VPWR u_rf.reg3_q\[20\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06640_ _01323_ _01860_ _01311_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_125_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
X_06571_ u_rf.reg12_q\[3\] _01608_ _01670_ u_rf.reg27_q\[3\] VGND VGND VPWR VPWR _01835_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_111_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08310_ u_rf.reg31_q\[7\] _03504_ _03505_ u_rf.reg11_q\[7\] _03506_ VGND VGND VPWR
+ VPWR _03507_ sky130_fd_sc_hd__a221o_1
X_09290_ _04385_ u_decod.rs2_data_q\[8\] _04386_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__and3_1
XFILLER_0_157_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_14 _01616_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08241_ u_rf.reg9_q\[4\] _03294_ _03296_ u_rf.reg20_q\[4\] VGND VGND VPWR VPWR _03441_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_36 _03274_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _02502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _03310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_31_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_69 _04409_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_83 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_58 _03366_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08172_ u_rf.reg6_q\[1\] _03304_ _03306_ u_rf.reg13_q\[1\] VGND VGND VPWR VPWR _03375_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07123_ u_rf.reg5_q\[14\] _01569_ _01556_ u_rf.reg6_q\[14\] VGND VGND VPWR VPWR _02365_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput110 net110 VGND VGND VPWR VPWR adr_o[18] sky130_fd_sc_hd__buf_2
X_07054_ net37 _02047_ _02049_ net54 _02051_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput121 net121 VGND VGND VPWR VPWR adr_o[28] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_140_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput143 net143 VGND VGND VPWR VPWR icache_adr_o[18] sky130_fd_sc_hd__buf_2
X_06005_ u_decod.rs2_data_q\[25\] u_decod.rs1_data_q\[25\] VGND VGND VPWR VPWR _01276_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput132 net132 VGND VGND VPWR VPWR adr_o[9] sky130_fd_sc_hd__buf_4
XFILLER_0_88_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput154 net154 VGND VGND VPWR VPWR icache_adr_o[28] sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_120_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput165 net165 VGND VGND VPWR VPWR icache_adr_o[9] sky130_fd_sc_hd__buf_4
Xoutput176 net176 VGND VGND VPWR VPWR store_data_o[18] sky130_fd_sc_hd__clkbuf_4
Xoutput187 net187 VGND VGND VPWR VPWR store_data_o[28] sky130_fd_sc_hd__buf_4
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput198 net198 VGND VGND VPWR VPWR store_data_o[9] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07956_ _02357_ u_decod.exe_ff_res_data_i\[31\] _03163_ VGND VGND VPWR VPWR _03164_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_145_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06907_ u_rf.reg6_q\[10\] _01554_ _01651_ u_rf.reg22_q\[10\] VGND VGND VPWR VPWR
+ _02157_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07887_ _02618_ _03097_ _02621_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09626_ u_rf.reg3_q\[17\] _04463_ _04582_ VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06838_ _01307_ _02059_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09557_ _04552_ VGND VGND VPWR VPWR _00081_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_65_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06769_ u_rf.reg26_q\[7\] _01640_ _01643_ u_rf.reg20_q\[7\] VGND VGND VPWR VPWR _02025_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_35_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09488_ _04515_ VGND VGND VPWR VPWR _00049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08508_ u_rf.reg30_q\[16\] _03281_ _03283_ u_rf.reg10_q\[16\] _03695_ VGND VGND VPWR
+ VPWR _03696_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08439_ u_rf.reg6_q\[13\] _03387_ _03270_ u_rf.reg8_q\[13\] _03629_ VGND VGND VPWR
+ VPWR _03630_ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11450_ _05592_ VGND VGND VPWR VPWR _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _05035_ VGND VGND VPWR VPWR _00442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11381_ u_rf.reg28_q\[6\] u_decod.rf_ff_res_data_i\[6\] _05549_ VGND VGND VPWR VPWR
+ _05556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10332_ u_decod.rf_ff_res_data_i\[28\] VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__buf_2
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12002_ clknet_leaf_83_clk u_exe.bu_pc_res\[15\] net366 VGND VGND VPWR VPWR u_exe.pc_data_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10263_ _04950_ VGND VGND VPWR VPWR _00389_ sky130_fd_sc_hd__clkbuf_1
X_10194_ _04740_ u_rf.reg11_q\[9\] _04900_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__mux2_1
Xfanout370 net371 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12904_ clknet_leaf_21_clk _00941_ net286 VGND VGND VPWR VPWR u_rf.reg29_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12835_ clknet_leaf_108_clk _00872_ net312 VGND VGND VPWR VPWR u_rf.reg27_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12766_ clknet_leaf_134_clk _00803_ net232 VGND VGND VPWR VPWR u_rf.reg25_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12697_ clknet_leaf_57_clk _00734_ net293 VGND VGND VPWR VPWR u_rf.reg22_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11717_ clknet_leaf_111_clk _00009_ net317 VGND VGND VPWR VPWR u_rf.reg2_q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11648_ u_decod.branch_imm_q_o\[3\] _01831_ _05696_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__mux2_1
Xinput12 icache_instr_i[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput34 load_data_i[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_1
Xinput45 load_data_i[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput23 icache_instr_i[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
X_11579_ _04728_ u_rf.reg31_q\[3\] _05657_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__mux2_1
Xinput78 reset_adr_i[21] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
Xinput89 reset_adr_i[31] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
XFILLER_0_107_492 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput67 reset_adr_i[11] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput56 load_data_i[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07810_ u_rf.reg7_q\[28\] _01562_ _01780_ u_rf.reg29_q\[28\] _03023_ VGND VGND VPWR
+ VPWR _03024_ sky130_fd_sc_hd__a221o_1
X_08790_ u_rf.reg6_q\[29\] _03304_ _03306_ u_rf.reg13_q\[29\] VGND VGND VPWR VPWR
+ _03965_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07741_ u_decod.pc_q_o\[27\] _02909_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07672_ u_rf.reg5_q\[25\] _01569_ _01606_ u_rf.reg3_q\[25\] _02891_ VGND VGND VPWR
+ VPWR _02892_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_140_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09411_ _04468_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__clkbuf_1
X_06623_ u_rf.reg23_q\[4\] _01613_ _01656_ u_rf.reg10_q\[4\] _01884_ VGND VGND VPWR
+ VPWR _01885_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_09342_ _04409_ u_decod.instr_operation_q\[0\] _04410_ VGND VGND VPWR VPWR _04420_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_59_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06554_ _01430_ _01259_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__nand2_2
XFILLER_0_118_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09273_ _04378_ _04381_ _04382_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06485_ u_decod.rs1_data_q\[9\] u_decod.rs1_data_q\[25\] _01702_ VGND VGND VPWR VPWR
+ _01752_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08224_ u_rf.reg27_q\[3\] _03365_ _03366_ u_rf.reg19_q\[3\] _03424_ VGND VGND VPWR
+ VPWR _03425_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08155_ u_rf.reg4_q\[1\] _03356_ _03357_ u_rf.reg17_q\[1\] VGND VGND VPWR VPWR _03358_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07106_ _01685_ _02137_ _02348_ _01458_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08086_ _03289_ VGND VGND VPWR VPWR _03290_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07037_ _02281_ _01347_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08988_ u_decod.rs1_data_q\[25\] u_decod.branch_imm_q_o\[25\] VGND VGND VPWR VPWR
+ _04138_ sky130_fd_sc_hd__nor2_1
X_07939_ u_rf.reg23_q\[31\] _02652_ _01654_ u_rf.reg22_q\[31\] _03146_ VGND VGND VPWR
+ VPWR _03147_ sky130_fd_sc_hd__a221o_1
X_10950_ _05327_ VGND VGND VPWR VPWR _00699_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10881_ _05290_ VGND VGND VPWR VPWR _00667_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ u_rf.reg3_q\[9\] _04446_ _04571_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__mux2_1
X_12620_ clknet_leaf_10_clk _00657_ net225 VGND VGND VPWR VPWR u_rf.reg20_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12551_ clknet_leaf_4_clk _00588_ net212 VGND VGND VPWR VPWR u_rf.reg18_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11502_ _05619_ VGND VGND VPWR VPWR _00959_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_198 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12482_ clknet_leaf_133_clk _00519_ net230 VGND VGND VPWR VPWR u_rf.reg16_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11433_ u_rf.reg28_q\[31\] u_decod.rf_ff_res_data_i\[31\] _05548_ VGND VGND VPWR
+ VPWR _05583_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_541 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_78_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11364_ _05546_ VGND VGND VPWR VPWR _00894_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10315_ u_rf.reg12_q\[22\] _04985_ _04981_ VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__mux2_1
X_11295_ u_rf.reg26_q\[30\] u_decod.rf_ff_res_data_i\[30\] _05476_ VGND VGND VPWR
+ VPWR _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_257 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_109_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10177_ _04901_ VGND VGND VPWR VPWR _00352_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_471 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12818_ clknet_leaf_41_clk _00855_ net278 VGND VGND VPWR VPWR u_rf.reg26_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12749_ clknet_leaf_5_clk _00786_ net216 VGND VGND VPWR VPWR u_rf.reg24_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_340 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06270_ _01536_ _01537_ _01538_ _01539_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_213 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09960_ _04783_ VGND VGND VPWR VPWR _00253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08911_ _01292_ u_decod.branch_imm_q_o\[14\] VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__or2_1
X_09891_ _04736_ u_rf.reg7_q\[7\] _04722_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__mux2_1
X_08842_ u_decod.rs1_data_q\[4\] u_decod.branch_imm_q_o\[4\] VGND VGND VPWR VPWR _04013_
+ sky130_fd_sc_hd__nand2_1
X_08773_ u_rf.reg16_q\[28\] _03322_ _03515_ u_rf.reg5_q\[28\] VGND VGND VPWR VPWR
+ _03949_ sky130_fd_sc_hd__a22o_1
X_05985_ u_decod.rd_v_q _01056_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__nand2_1
X_07724_ u_rf.reg30_q\[26\] _01581_ _02419_ u_rf.reg28_q\[26\] VGND VGND VPWR VPWR
+ _02942_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_706 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07655_ _02835_ _02875_ _02189_ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06606_ _01449_ _01868_ _01464_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07586_ _02803_ _02805_ _02807_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09325_ _04411_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_90_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06537_ _01737_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_157_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09256_ _04368_ _04369_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06468_ _01726_ _01735_ _01679_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08207_ _03272_ VGND VGND VPWR VPWR _03408_ sky130_fd_sc_hd__buf_6
XFILLER_0_51_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_251 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09187_ _04100_ _04274_ _04275_ _04310_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[18\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06399_ _01538_ _01558_ _01573_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__and3_4
XFILLER_0_31_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08138_ _03280_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__buf_6
XFILLER_0_114_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_522 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08069_ _03272_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__buf_6
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11080_ _05396_ VGND VGND VPWR VPWR _00760_ sky130_fd_sc_hd__clkbuf_1
X_10100_ _04859_ VGND VGND VPWR VPWR _00317_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _04822_ VGND VGND VPWR VPWR _00285_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11982_ clknet_leaf_65_clk net436 net347 VGND VGND VPWR VPWR u_decod.pc_q_o\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_728 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10933_ _05318_ VGND VGND VPWR VPWR _00691_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10864_ _05281_ VGND VGND VPWR VPWR _00659_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10795_ u_rf.reg19_q\[19\] _04978_ _05235_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__mux2_1
X_12603_ clknet_leaf_122_clk _00640_ net241 VGND VGND VPWR VPWR u_rf.reg20_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12534_ clknet_leaf_48_clk _00571_ net300 VGND VGND VPWR VPWR u_rf.reg17_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12465_ clknet_leaf_54_clk _00502_ net296 VGND VGND VPWR VPWR u_rf.reg15_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11416_ _05574_ VGND VGND VPWR VPWR _00918_ sky130_fd_sc_hd__clkbuf_1
X_12396_ clknet_leaf_10_clk _00433_ net225 VGND VGND VPWR VPWR u_rf.reg13_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11347_ _04768_ u_rf.reg27_q\[22\] _05535_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11278_ _05501_ VGND VGND VPWR VPWR _00853_ sky130_fd_sc_hd__clkbuf_1
X_13017_ clknet_leaf_65_clk _01054_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[30\]
+ sky130_fd_sc_hd__dfxtp_1
X_10229_ _04928_ VGND VGND VPWR VPWR _00377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05770_ u_decod.dec0.instr_i\[0\] u_decod.dec0.funct3\[2\] VGND VGND VPWR VPWR _01093_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_77_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07440_ u_decod.rf_ff_res_data_i\[20\] _01550_ _01773_ _02647_ _02669_ VGND VGND
+ VPWR VPWR _02670_ sky130_fd_sc_hd__a221o_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07371_ _02596_ _02598_ _02600_ _02602_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__or4_1
X_09110_ u_decod.pc_q_o\[8\] u_decod.branch_imm_q_o\[8\] VGND VGND VPWR VPWR _04244_
+ sky130_fd_sc_hd__or2_1
X_06322_ _01591_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_40_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_896 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09041_ _01266_ _01273_ _01277_ _01286_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06253_ u_decod.dec0.instr_i\[21\] _01521_ u_decod.exe_ff_rd_adr_q_i\[2\] _01522_
+ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06184_ u_decod.rs2_data_q\[3\] VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_352 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09943_ u_decod.rf_ff_res_data_i\[24\] VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09874_ _04725_ VGND VGND VPWR VPWR _00225_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08825_ _02621_ VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_51_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _03926_ _03928_ _03930_ _03932_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__or4_1
X_05968_ _01079_ _01220_ _01245_ _01234_ VGND VGND VPWR VPWR u_decod.dec0.operation_o\[2\]
+ sky130_fd_sc_hd__a22o_1
X_08687_ u_rf.reg16_q\[24\] _03322_ _03324_ u_rf.reg5_q\[24\] VGND VGND VPWR VPWR
+ _03867_ sky130_fd_sc_hd__a22o_1
X_05899_ net506 _01118_ _01119_ net86 _01191_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__a221o_1
X_07707_ _02618_ _02925_ _02621_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__a21oi_1
X_07638_ _02850_ _02859_ _02359_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__o21a_1
X_07569_ u_rf.reg30_q\[23\] _01581_ _02419_ u_rf.reg28_q\[23\] VGND VGND VPWR VPWR
+ _02793_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09308_ _04397_ u_decod.rs2_data_q\[16\] _04398_ VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__and3_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10580_ _05131_ VGND VGND VPWR VPWR _00525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09239_ _04146_ _04206_ _04197_ _04354_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[26\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12250_ clknet_leaf_60_clk _00287_ net340 VGND VGND VPWR VPWR u_rf.reg8_q\[31\] sky130_fd_sc_hd__dfrtp_1
X_12181_ clknet_leaf_46_clk _00218_ net298 VGND VGND VPWR VPWR u_rf.reg6_q\[26\] sky130_fd_sc_hd__dfrtp_1
X_11201_ _05460_ VGND VGND VPWR VPWR _00817_ sky130_fd_sc_hd__clkbuf_1
X_11132_ u_rf.reg24_q\[17\] _04974_ _05416_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11063_ _05387_ VGND VGND VPWR VPWR _00752_ sky130_fd_sc_hd__clkbuf_1
X_10014_ u_rf.reg8_q\[21\] _04472_ _04812_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11965_ clknet_leaf_84_clk net444 net366 VGND VGND VPWR VPWR u_decod.pc_q_o\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_739 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10916_ u_rf.reg21_q\[11\] _04962_ _05308_ VGND VGND VPWR VPWR _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11896_ clknet_leaf_96_clk u_decod.rs2_data_nxt\[17\] net332 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10847_ u_rf.reg20_q\[11\] _04962_ _05271_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10778_ _05236_ VGND VGND VPWR VPWR _00618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12517_ clknet_leaf_124_clk _00554_ net239 VGND VGND VPWR VPWR u_rf.reg17_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12448_ clknet_leaf_115_clk _00485_ net324 VGND VGND VPWR VPWR u_rf.reg15_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ clknet_leaf_11_clk _00416_ net222 VGND VGND VPWR VPWR u_rf.reg13_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06940_ _01479_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06871_ u_rf.reg7_q\[9\] _01559_ _01604_ u_rf.reg3_q\[9\] VGND VGND VPWR VPWR _02123_
+ sky130_fd_sc_hd__a22o_1
X_08610_ _03178_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__clkbuf_4
X_05822_ u_decod.pc0_q_i\[11\] _01129_ VGND VGND VPWR VPWR _01133_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09590_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__buf_6
X_08541_ _03721_ _03723_ _03725_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__or4_1
X_05753_ u_decod.dec0.funct3\[1\] VGND VGND VPWR VPWR _01076_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08472_ u_rf.reg15_q\[14\] _03300_ _03302_ u_rf.reg24_q\[14\] _03661_ VGND VGND VPWR
+ VPWR _03662_ sky130_fd_sc_hd__a221o_1
X_07423_ u_rf.reg6_q\[20\] _01556_ _01584_ u_rf.reg11_q\[20\] VGND VGND VPWR VPWR
+ _02653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_324 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_302 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07354_ _01423_ _02585_ _02586_ _01505_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07285_ u_rf.reg23_q\[17\] _01612_ _01621_ u_rf.reg24_q\[17\] VGND VGND VPWR VPWR
+ _02521_ sky130_fd_sc_hd__a22o_1
X_06305_ _01574_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__buf_6
XFILLER_0_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09024_ _04161_ _04164_ _04162_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_103_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06236_ _01424_ _01496_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06167_ _01435_ _01437_ _01314_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06098_ u_decod.rs2_data_q\[23\] _01367_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09926_ _04760_ VGND VGND VPWR VPWR _00242_ sky130_fd_sc_hd__clkbuf_1
X_09857_ _04714_ VGND VGND VPWR VPWR _00219_ sky130_fd_sc_hd__clkbuf_1
X_09788_ _04677_ VGND VGND VPWR VPWR _00187_ sky130_fd_sc_hd__clkbuf_1
X_08808_ u_rf.reg18_q\[30\] _03352_ _03354_ u_rf.reg23_q\[30\] _03981_ VGND VGND VPWR
+ VPWR _03982_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ u_rf.reg22_q\[27\] _03274_ _03410_ u_rf.reg3_q\[27\] VGND VGND VPWR VPWR
+ _03916_ sky130_fd_sc_hd__a22o_1
XANTENNA_104 u_decod.dec0.funct7\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_115 u_decod.rs1_data_q\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _01780_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 _03310_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 _01384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ clknet_leaf_122_clk _00042_ net247 VGND VGND VPWR VPWR u_rf.reg1_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10701_ _05195_ VGND VGND VPWR VPWR _00582_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_159 _05632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11681_ u_decod.branch_imm_q_o\[19\] _02594_ _05696_ VGND VGND VPWR VPWR _05715_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ u_rf.reg17_q\[6\] _04951_ _05152_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10563_ _05122_ VGND VGND VPWR VPWR _00517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12302_ clknet_leaf_6_clk _00339_ net216 VGND VGND VPWR VPWR u_rf.reg10_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10494_ _04734_ u_rf.reg15_q\[6\] _05078_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12233_ clknet_leaf_24_clk _00270_ net266 VGND VGND VPWR VPWR u_rf.reg8_q\[14\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_15_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12164_ clknet_leaf_106_clk _00201_ net319 VGND VGND VPWR VPWR u_rf.reg6_q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ clknet_leaf_137_clk _00132_ net206 VGND VGND VPWR VPWR u_rf.reg4_q\[4\] sky130_fd_sc_hd__dfrtp_1
X_11115_ u_rf.reg24_q\[9\] _04957_ _05405_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__mux2_1
X_11046_ _05378_ VGND VGND VPWR VPWR _00744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12997_ clknet_leaf_92_clk _01034_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[10\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_424 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11948_ clknet_leaf_95_clk u_decod.dec0.rd_o\[2\] net325 VGND VGND VPWR VPWR u_decod.exe_ff_rd_adr_q_i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_156_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11879_ clknet_leaf_99_clk u_decod.rs2_data_nxt\[0\] net329 VGND VGND VPWR VPWR u_decod.rs2_data_q\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07070_ u_rf.reg19_q\[13\] _01594_ _01649_ u_rf.reg4_q\[13\] VGND VGND VPWR VPWR
+ _02314_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_611 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06021_ u_decod.rs1_data_q\[14\] VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09711_ _04635_ VGND VGND VPWR VPWR _00152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07972_ _01204_ _01226_ _03169_ _03177_ VGND VGND VPWR VPWR _03178_ sky130_fd_sc_hd__o31a_4
X_06923_ u_rf.reg25_q\[10\] _01574_ _01620_ u_rf.reg24_q\[10\] _02172_ VGND VGND VPWR
+ VPWR _02173_ sky130_fd_sc_hd__a221o_1
X_09642_ _04598_ VGND VGND VPWR VPWR _00120_ sky130_fd_sc_hd__clkbuf_1
X_06854_ _01305_ _01428_ _01434_ _01337_ _02106_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__a221oi_2
X_09573_ net530 _04480_ _04555_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__mux2_1
X_05805_ _01099_ _01116_ _01117_ _01120_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__a31o_2
X_06785_ _01951_ _02039_ _01315_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_143_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05736_ u_decod.branch_imm_q_o\[0\] _01061_ VGND VGND VPWR VPWR _01062_ sky130_fd_sc_hd__nand2_1
X_08524_ u_rf.reg26_q\[17\] _03344_ _03345_ u_rf.reg21_q\[17\] VGND VGND VPWR VPWR
+ _03711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08455_ u_decod.rf_ff_res_data_i\[13\] _03382_ _03645_ _03404_ VGND VGND VPWR VPWR
+ _03646_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07406_ _01405_ _02635_ _01366_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_63_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_742 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08386_ u_rf.reg27_q\[10\] _03319_ _03321_ u_rf.reg19_q\[10\] _03579_ VGND VGND VPWR
+ VPWR _03580_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07337_ u_decod.rf_ff_res_data_i\[18\] _01550_ _01773_ _02551_ _02570_ VGND VGND
+ VPWR VPWR _02571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_847 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07268_ _01059_ _02492_ _02497_ _02504_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09007_ _04142_ _04148_ _04147_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_104_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07199_ u_decod.rf_ff_res_data_i\[15\] _01550_ u_decod.exe_ff_res_data_i\[15\] _01772_
+ _02438_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__a221o_1
X_06219_ net98 _01063_ net101 VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09909_ u_decod.rf_ff_res_data_i\[13\] VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__buf_2
X_12920_ clknet_leaf_67_clk _00957_ net349 VGND VGND VPWR VPWR u_rf.reg29_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_12851_ clknet_leaf_68_clk _00888_ net351 VGND VGND VPWR VPWR u_rf.reg27_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_11802_ clknet_leaf_81_clk net155 net368 VGND VGND VPWR VPWR u_decod.pc0_q_i\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ clknet_leaf_28_clk _00819_ net257 VGND VGND VPWR VPWR u_rf.reg25_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11733_ clknet_leaf_32_clk _00025_ net262 VGND VGND VPWR VPWR u_rf.reg2_q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11664_ _01079_ _05700_ _02644_ _05706_ VGND VGND VPWR VPWR _01034_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10615_ _05149_ VGND VGND VPWR VPWR _00542_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11595_ _05669_ VGND VGND VPWR VPWR _01002_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10546_ _04786_ u_rf.reg15_q\[31\] _05077_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10477_ _05075_ VGND VGND VPWR VPWR _00478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12216_ clknet_leaf_57_clk _00253_ net292 VGND VGND VPWR VPWR u_rf.reg7_q\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12147_ clknet_leaf_66_clk _00184_ net356 VGND VGND VPWR VPWR u_rf.reg5_q\[24\] sky130_fd_sc_hd__dfrtp_1
X_12078_ clknet_leaf_28_clk _00115_ net256 VGND VGND VPWR VPWR u_rf.reg3_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11029_ _04719_ u_rf.reg23_q\[0\] _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06570_ u_rf.reg16_q\[3\] _01564_ _01592_ u_rf.reg18_q\[3\] _01833_ VGND VGND VPWR
+ VPWR _01834_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08240_ u_rf.reg30_q\[4\] _03281_ _03283_ u_rf.reg10_q\[4\] _03439_ VGND VGND VPWR
+ VPWR _03440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_37 _03276_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_48 _03311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _01630_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08171_ _03302_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__buf_8
XANTENNA_26 _03176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07122_ _01639_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_59 _03373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_113_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_95 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07053_ _01422_ _02296_ _02297_ _01505_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR access_size_o[2] sky130_fd_sc_hd__buf_4
XFILLER_0_31_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 net122 VGND VGND VPWR VPWR adr_o[29] sky130_fd_sc_hd__buf_4
Xoutput111 net111 VGND VGND VPWR VPWR adr_o[19] sky130_fd_sc_hd__buf_2
X_06004_ u_decod.rs2_data_q\[25\] u_decod.rs1_data_q\[25\] VGND VGND VPWR VPWR _01275_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_88_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput133 net133 VGND VGND VPWR VPWR adr_v_o sky130_fd_sc_hd__buf_4
Xoutput144 net144 VGND VGND VPWR VPWR icache_adr_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_140_496 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput155 net155 VGND VGND VPWR VPWR icache_adr_o[29] sky130_fd_sc_hd__buf_2
Xoutput166 net166 VGND VGND VPWR VPWR is_store_o sky130_fd_sc_hd__buf_2
XFILLER_0_56_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput177 net177 VGND VGND VPWR VPWR store_data_o[19] sky130_fd_sc_hd__buf_4
XFILLER_0_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput188 net188 VGND VGND VPWR VPWR store_data_o[29] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_145_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07955_ u_decod.rf_ff_res_data_i\[31\] _02358_ _02743_ _03143_ _03162_ VGND VGND
+ VPWR VPWR _03163_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_145_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06906_ _02156_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[10\] sky130_fd_sc_hd__inv_2
X_07886_ _02619_ net56 VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09625_ _04589_ VGND VGND VPWR VPWR _00112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06837_ _02084_ _02090_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[8\] sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09556_ u_rf.reg0_q\[17\] _04463_ _04544_ VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06768_ u_rf.reg15_q\[7\] _01600_ _01670_ u_rf.reg27_q\[7\] _02023_ VGND VGND VPWR
+ VPWR _02024_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09487_ u_rf.reg1_q\[17\] _04463_ _04507_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__mux2_1
X_06699_ _01825_ _01866_ _01906_ _01957_ _01479_ _01476_ VGND VGND VPWR VPWR _01958_
+ sky130_fd_sc_hd__mux4_1
X_08507_ u_rf.reg26_q\[16\] _03343_ _03286_ u_rf.reg21_q\[16\] VGND VGND VPWR VPWR
+ _03695_ sky130_fd_sc_hd__a22o_1
X_08438_ u_rf.reg27_q\[13\] _03246_ _03247_ u_rf.reg19_q\[13\] VGND VGND VPWR VPWR
+ _03629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08369_ u_decod.exe_ff_res_data_i\[9\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[9\]
+ _03563_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a221o_1
X_10400_ _04776_ u_rf.reg13_q\[26\] _05028_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11380_ _05555_ VGND VGND VPWR VPWR _00901_ sky130_fd_sc_hd__clkbuf_1
X_10331_ _04996_ VGND VGND VPWR VPWR _00411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10262_ u_rf.reg12_q\[5\] _04949_ _04939_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__mux2_1
X_12001_ clknet_leaf_82_clk u_exe.bu_pc_res\[14\] net366 VGND VGND VPWR VPWR u_exe.pc_data_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10193_ _04909_ VGND VGND VPWR VPWR _00360_ sky130_fd_sc_hd__clkbuf_1
Xfanout371 net372 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12903_ clknet_leaf_3_clk _00940_ net213 VGND VGND VPWR VPWR u_rf.reg29_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_12834_ clknet_leaf_130_clk _00871_ net230 VGND VGND VPWR VPWR u_rf.reg27_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12765_ clknet_leaf_15_clk _00802_ net281 VGND VGND VPWR VPWR u_rf.reg25_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11716_ clknet_leaf_107_clk _00008_ net314 VGND VGND VPWR VPWR u_rf.reg2_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12696_ clknet_leaf_62_clk _00733_ net343 VGND VGND VPWR VPWR u_rf.reg22_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11647_ _05697_ VGND VGND VPWR VPWR _01026_ sky130_fd_sc_hd__clkbuf_1
Xinput13 icache_instr_i[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
XFILLER_0_107_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _05660_ VGND VGND VPWR VPWR _00994_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput35 load_data_i[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput24 icache_instr_i[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
Xinput46 load_data_i[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput79 reset_adr_i[22] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
X_10529_ _05103_ VGND VGND VPWR VPWR _00502_ sky130_fd_sc_hd__clkbuf_1
Xinput68 reset_adr_i[12] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput57 load_data_i[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_2
XFILLER_0_149_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_856 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07740_ u_decod.pc_q_o\[27\] _02909_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__or2_1
X_07671_ u_rf.reg15_q\[25\] _01600_ _01612_ u_rf.reg23_q\[25\] VGND VGND VPWR VPWR
+ _02891_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09410_ u_rf.reg2_q\[19\] _04467_ _04449_ VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__mux2_1
X_06622_ u_rf.reg6_q\[4\] _01555_ _01652_ u_rf.reg22_q\[4\] VGND VGND VPWR VPWR _01884_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09341_ _04419_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlymetal6s2s_1
X_06553_ _01484_ _01816_ _01817_ _01813_ _01435_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__a32o_1
XFILLER_0_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09272_ _04378_ _04381_ _04382_ VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__nand3_1
XFILLER_0_114_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06484_ _01747_ _01501_ _01706_ _01750_ _01480_ _01477_ VGND VGND VPWR VPWR _01751_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_466 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08223_ u_rf.reg16_q\[3\] _03322_ _03324_ u_rf.reg5_q\[3\] VGND VGND VPWR VPWR _03424_
+ sky130_fd_sc_hd__a22o_1
X_08154_ _03266_ VGND VGND VPWR VPWR _03357_ sky130_fd_sc_hd__buf_12
XTAP_TAPCELL_ROW_155_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08085_ _03210_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__clkbuf_8
X_07105_ _01455_ _01754_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07036_ _01298_ _02231_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_58_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08987_ u_decod.rs1_data_q\[25\] u_decod.branch_imm_q_o\[25\] VGND VGND VPWR VPWR
+ _04137_ sky130_fd_sc_hd__and2_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ u_rf.reg6_q\[31\] _01557_ _02375_ u_rf.reg11_q\[31\] VGND VGND VPWR VPWR
+ _03146_ sky130_fd_sc_hd__a22o_1
X_07869_ _02357_ u_decod.exe_ff_res_data_i\[29\] _03080_ VGND VGND VPWR VPWR _03081_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_97_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10880_ u_rf.reg20_q\[27\] _04995_ _05282_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__mux2_1
X_09608_ _04580_ VGND VGND VPWR VPWR _00104_ sky130_fd_sc_hd__clkbuf_1
X_09539_ u_rf.reg0_q\[9\] _04446_ _04533_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12550_ clknet_leaf_139_clk _00587_ net203 VGND VGND VPWR VPWR u_rf.reg18_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11501_ _04786_ u_rf.reg29_q\[31\] _05584_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__mux2_1
X_12481_ clknet_leaf_118_clk _00518_ net326 VGND VGND VPWR VPWR u_rf.reg16_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_514 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11432_ _05582_ VGND VGND VPWR VPWR _00926_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_203 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11363_ _04784_ u_rf.reg27_q\[30\] _05512_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11294_ _05509_ VGND VGND VPWR VPWR _00861_ sky130_fd_sc_hd__clkbuf_1
X_10314_ u_decod.rf_ff_res_data_i\[22\] VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__buf_2
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10245_ _04423_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__nor2_4
X_10176_ _04719_ u_rf.reg11_q\[0\] _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_704 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12817_ clknet_leaf_57_clk _00854_ net293 VGND VGND VPWR VPWR u_rf.reg26_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12748_ clknet_leaf_25_clk _00785_ net265 VGND VGND VPWR VPWR u_rf.reg24_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_648 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_328 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12679_ clknet_leaf_3_clk _00716_ net213 VGND VGND VPWR VPWR u_rf.reg22_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_136 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08910_ _04042_ _04071_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__nor2_1
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09890_ u_decod.rf_ff_res_data_i\[7\] VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08841_ u_decod.rs1_data_q\[4\] u_decod.branch_imm_q_o\[4\] VGND VGND VPWR VPWR _04012_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_76 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08772_ u_rf.reg7_q\[28\] _03369_ _03370_ u_rf.reg25_q\[28\] _03947_ VGND VGND VPWR
+ VPWR _03948_ sky130_fd_sc_hd__a221o_1
X_05984_ _01256_ VGND VGND VPWR VPWR u_decod.dec0.access_size_o\[2\] sky130_fd_sc_hd__clkbuf_1
X_07723_ u_rf.reg17_q\[26\] _02379_ _02360_ u_rf.reg9_q\[26\] _02940_ VGND VGND VPWR
+ VPWR _02941_ sky130_fd_sc_hd__a221o_1
X_07654_ _02584_ _02684_ _02778_ _02874_ _01475_ _02685_ VGND VGND VPWR VPWR _02875_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06605_ u_decod.rs1_data_q\[19\] _01683_ u_decod.rs1_data_q\[11\] u_decod.rs1_data_q\[27\]
+ _01702_ _01684_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__mux4_1
X_07585_ u_rf.reg29_q\[23\] _01780_ _02364_ u_rf.reg21_q\[23\] _02808_ VGND VGND VPWR
+ VPWR _02809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09324_ _04409_ u_decod.rs2_data_q\[23\] _04410_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__and3_1
X_06536_ _01772_ u_decod.exe_ff_res_data_i\[2\] _01775_ _01801_ VGND VGND VPWR VPWR
+ _01802_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09255_ u_decod.pc_q_o\[28\] u_decod.branch_imm_q_o\[28\] VGND VGND VPWR VPWR _04369_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06467_ _01728_ _01730_ _01732_ _01734_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__or4_1
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08206_ _03270_ VGND VGND VPWR VPWR _03407_ sky130_fd_sc_hd__buf_8
XFILLER_0_7_263 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09186_ _04308_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__xor2_1
X_06398_ _01667_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__buf_8
XFILLER_0_44_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08137_ u_decod.pc0_q_i\[0\] _03259_ _03339_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[0\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_534 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08068_ _03217_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__buf_6
XFILLER_0_101_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07019_ u_rf.reg3_q\[12\] _01606_ _01639_ u_rf.reg21_q\[12\] _02264_ VGND VGND VPWR
+ VPWR _02265_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10030_ u_rf.reg8_q\[29\] _04488_ _04812_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ clknet_leaf_65_clk net435 net357 VGND VGND VPWR VPWR u_decod.pc_q_o\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ u_rf.reg21_q\[19\] _04978_ _05308_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10863_ u_rf.reg20_q\[19\] _04978_ _05271_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ clknet_leaf_59_clk _00639_ net292 VGND VGND VPWR VPWR u_rf.reg19_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_762 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10794_ _05244_ VGND VGND VPWR VPWR _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12533_ clknet_leaf_44_clk _00570_ net295 VGND VGND VPWR VPWR u_rf.reg17_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12464_ clknet_leaf_36_clk _00501_ net273 VGND VGND VPWR VPWR u_rf.reg15_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11415_ u_rf.reg28_q\[22\] u_decod.rf_ff_res_data_i\[22\] _05571_ VGND VGND VPWR
+ VPWR _05574_ sky130_fd_sc_hd__mux2_1
X_12395_ clknet_leaf_135_clk _00432_ net207 VGND VGND VPWR VPWR u_rf.reg13_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11346_ _05537_ VGND VGND VPWR VPWR _00885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13016_ clknet_leaf_65_clk _01053_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[29\]
+ sky130_fd_sc_hd__dfxtp_1
X_11277_ u_rf.reg26_q\[21\] u_decod.rf_ff_res_data_i\[21\] _05499_ VGND VGND VPWR
+ VPWR _05501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10228_ _04774_ u_rf.reg11_q\[25\] _04922_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__mux2_1
X_10159_ u_rf.reg10_q\[25\] _04480_ _04885_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_420 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07370_ u_rf.reg5_q\[19\] _01569_ _01562_ u_rf.reg7_q\[19\] _02601_ VGND VGND VPWR
+ VPWR _02602_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06321_ _01590_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__buf_6
XFILLER_0_127_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09040_ _04179_ _04180_ _04181_ _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06252_ u_decod.dec0.instr_i\[22\] VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06183_ _01445_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09942_ _04771_ VGND VGND VPWR VPWR _00247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _04724_ u_rf.reg7_q\[1\] _04722_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__mux2_1
X_08824_ net435 _03257_ _03997_ _03178_ VGND VGND VPWR VPWR u_decod.rs1_data\[30\]
+ sky130_fd_sc_hd__a22o_1
X_08755_ u_rf.reg0_q\[27\] _03420_ _03421_ u_rf.reg12_q\[27\] _03931_ VGND VGND VPWR
+ VPWR _03932_ sky130_fd_sc_hd__a221o_1
X_07706_ _02619_ net51 VGND VGND VPWR VPWR _02925_ sky130_fd_sc_hd__nand2_1
X_05967_ _01075_ _01084_ _01091_ _01243_ _01244_ VGND VGND VPWR VPWR _01245_ sky130_fd_sc_hd__a311o_1
X_08686_ u_rf.reg0_q\[24\] _03175_ _03328_ u_rf.reg12_q\[24\] _03865_ VGND VGND VPWR
+ VPWR _03866_ sky130_fd_sc_hd__a221o_1
X_05898_ _01189_ _01190_ VGND VGND VPWR VPWR _01191_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07637_ _02852_ _02854_ _02856_ _02858_ VGND VGND VPWR VPWR _02859_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07568_ u_decod.dec0.instr_i\[23\] _01206_ _02646_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_24_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09307_ _04401_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
X_06519_ u_rf.reg26_q\[2\] _01642_ _01645_ u_rf.reg20_q\[2\] VGND VGND VPWR VPWR _01785_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07499_ _01469_ _02137_ _01498_ _01905_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__o211a_1
X_09238_ _04352_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09169_ u_decod.pc_q_o\[16\] u_decod.branch_imm_q_o\[16\] VGND VGND VPWR VPWR _04295_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12180_ clknet_leaf_32_clk _00217_ net262 VGND VGND VPWR VPWR u_rf.reg6_q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11200_ u_rf.reg25_q\[17\] _04974_ _05452_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__mux2_1
X_11131_ _05423_ VGND VGND VPWR VPWR _00784_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_79_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11062_ _04755_ u_rf.reg23_q\[16\] _05380_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__mux2_1
X_10013_ _04813_ VGND VGND VPWR VPWR _00276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11964_ clknet_leaf_82_clk net450 net366 VGND VGND VPWR VPWR u_decod.pc_q_o\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11895_ clknet_leaf_97_clk u_decod.rs2_data_nxt\[16\] net332 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10915_ _05309_ VGND VGND VPWR VPWR _00682_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_88_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10846_ _05272_ VGND VGND VPWR VPWR _00650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_650 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10777_ u_rf.reg19_q\[10\] _04959_ _05235_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12516_ clknet_leaf_112_clk _00553_ net317 VGND VGND VPWR VPWR u_rf.reg17_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_117_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12447_ clknet_leaf_137_clk _00484_ net206 VGND VGND VPWR VPWR u_rf.reg15_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12378_ clknet_leaf_59_clk _00415_ net340 VGND VGND VPWR VPWR u_rf.reg12_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11329_ _05528_ VGND VGND VPWR VPWR _00877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_548 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06870_ u_rf.reg5_q\[9\] _01567_ _01593_ u_rf.reg19_q\[9\] _02121_ VGND VGND VPWR
+ VPWR _02122_ sky130_fd_sc_hd__a221o_1
X_05821_ _01100_ VGND VGND VPWR VPWR _01132_ sky130_fd_sc_hd__clkbuf_4
X_08540_ u_rf.reg27_q\[17\] _03318_ _03320_ u_rf.reg19_q\[17\] _03726_ VGND VGND VPWR
+ VPWR _03727_ sky130_fd_sc_hd__a221o_1
X_05752_ u_decod.dec0.instr_i\[4\] u_decod.dec0.instr_i\[5\] _01074_ VGND VGND VPWR
+ VPWR _01075_ sky130_fd_sc_hd__and3_2
X_08471_ u_rf.reg6_q\[14\] _03235_ _03236_ u_rf.reg13_q\[14\] VGND VGND VPWR VPWR
+ _03661_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07422_ _01613_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07353_ _01423_ _02543_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_300 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07284_ _02513_ _02515_ _02517_ _02519_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06304_ _01572_ _01566_ _01573_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_150_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09023_ _04166_ _04167_ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06235_ _01505_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_143_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06166_ _01436_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06097_ u_decod.rs2_data_q\[23\] _01367_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_53_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09925_ _04759_ u_rf.reg7_q\[18\] _04743_ VGND VGND VPWR VPWR _04760_ sky130_fd_sc_hd__mux2_1
X_09856_ u_rf.reg6_q\[27\] _04484_ _04706_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__mux2_1
X_08807_ u_rf.reg4_q\[30\] _03264_ _03266_ u_rf.reg17_q\[30\] VGND VGND VPWR VPWR
+ _03981_ sky130_fd_sc_hd__a22o_1
X_09787_ u_rf.reg5_q\[27\] _04484_ _04669_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__mux2_1
X_06999_ _01820_ _02245_ _01349_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ net464 _03773_ _03915_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[26\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_116 u_rf.reg0_q\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_105 u_decod.pc0_q_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 _01787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08669_ u_rf.reg27_q\[23\] _03365_ _03366_ u_rf.reg19_q\[23\] _03849_ VGND VGND VPWR
+ VPWR _03850_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 _01384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 _03331_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ u_rf.reg18_q\[6\] _04951_ _05188_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11680_ _05714_ VGND VGND VPWR VPWR _01042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_592 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10631_ _05158_ VGND VGND VPWR VPWR _00549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10562_ u_rf.reg16_q\[5\] _04949_ _05116_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__mux2_1
X_12301_ clknet_leaf_6_clk _00338_ net216 VGND VGND VPWR VPWR u_rf.reg10_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12232_ clknet_leaf_19_clk _00269_ net281 VGND VGND VPWR VPWR u_rf.reg8_q\[13\] sky130_fd_sc_hd__dfrtp_1
X_10493_ _05084_ VGND VGND VPWR VPWR _00485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12163_ clknet_leaf_107_clk _00200_ net319 VGND VGND VPWR VPWR u_rf.reg6_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_892 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _05414_ VGND VGND VPWR VPWR _00776_ sky130_fd_sc_hd__clkbuf_1
X_12094_ clknet_leaf_134_clk _00131_ net209 VGND VGND VPWR VPWR u_rf.reg4_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_11045_ _04738_ u_rf.reg23_q\[8\] _05369_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12996_ clknet_leaf_92_clk _01033_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[9\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11947_ clknet_leaf_95_clk u_decod.dec0.rd_o\[1\] net331 VGND VGND VPWR VPWR u_decod.exe_ff_rd_adr_q_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11878_ clknet_leaf_103_clk u_decod.dec0.access_size_o\[2\] net335 VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10829_ _05263_ VGND VGND VPWR VPWR _00642_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_491 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_478 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_623 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06020_ u_decod.rs2_data_q\[15\] _01289_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07971_ _03176_ VGND VGND VPWR VPWR _03177_ sky130_fd_sc_hd__inv_2
X_09710_ u_rf.reg4_q\[24\] _04478_ _04630_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__mux2_1
X_06922_ u_rf.reg26_q\[10\] _01640_ _01643_ u_rf.reg20_q\[10\] VGND VGND VPWR VPWR
+ _02172_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_147_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ net528 _04478_ _04593_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__mux2_1
X_06853_ _01306_ _01819_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__nor2_1
X_09572_ _04560_ VGND VGND VPWR VPWR _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05804_ u_exe.pc_data_q\[6\] _01118_ _01119_ net93 VGND VGND VPWR VPWR _01120_ sky130_fd_sc_hd__a22o_1
X_06784_ _01868_ _02038_ _01450_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ u_decod.pc0_q_i\[16\] _03565_ _03710_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[16\]
+ sky130_fd_sc_hd__a22o_1
X_05735_ u_decod.rs1_data_q\[0\] VGND VGND VPWR VPWR _01061_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08454_ _03635_ _03644_ VGND VGND VPWR VPWR _03645_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07405_ _01366_ _01405_ _02635_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08385_ u_rf.reg16_q\[10\] _03450_ _03515_ u_rf.reg5_q\[10\] VGND VGND VPWR VPWR
+ _03579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07336_ _02560_ _02569_ _01680_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_63_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_456 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09006_ u_decod.rs1_data_q\[24\] u_decod.branch_imm_q_o\[24\] _04137_ VGND VGND VPWR
+ VPWR _04153_ sky130_fd_sc_hd__a21oi_1
X_07267_ u_decod.rs2_data_q\[17\] _01380_ _01429_ _02502_ _02503_ VGND VGND VPWR VPWR
+ _02504_ sky130_fd_sc_hd__a311o_1
XFILLER_0_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07198_ _02421_ _02428_ _02437_ _01680_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__o31a_2
X_06218_ _01063_ net101 net98 VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__and3b_2
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06149_ _01394_ _01408_ _01418_ _01419_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__a31o_1
X_09908_ _04748_ VGND VGND VPWR VPWR _00236_ sky130_fd_sc_hd__clkbuf_1
X_09839_ u_rf.reg6_q\[19\] _04467_ _04695_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
X_12850_ clknet_leaf_39_clk _00887_ net279 VGND VGND VPWR VPWR u_rf.reg27_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11801_ clknet_leaf_76_clk net154 net368 VGND VGND VPWR VPWR u_decod.pc0_q_i\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ clknet_leaf_5_clk _00818_ net217 VGND VGND VPWR VPWR u_rf.reg25_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_11732_ clknet_leaf_67_clk _00024_ net349 VGND VGND VPWR VPWR u_rf.reg2_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11663_ _05693_ u_decod.branch_imm_q_o\[10\] VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__and2b_1
XFILLER_0_154_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10614_ u_rf.reg16_q\[30\] _05001_ _05115_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _04742_ u_rf.reg31_q\[10\] _05668_ VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10545_ _05111_ VGND VGND VPWR VPWR _00510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_130_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_130_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10476_ _04784_ u_rf.reg14_q\[30\] _05041_ VGND VGND VPWR VPWR _05075_ sky130_fd_sc_hd__mux2_1
X_12215_ clknet_leaf_71_clk _00252_ net353 VGND VGND VPWR VPWR u_rf.reg7_q\[28\] sky130_fd_sc_hd__dfrtp_1
X_12146_ clknet_leaf_38_clk _00183_ net277 VGND VGND VPWR VPWR u_rf.reg5_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12077_ clknet_leaf_5_clk _00114_ net215 VGND VGND VPWR VPWR u_rf.reg3_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11028_ _05368_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12979_ clknet_leaf_51_clk _01016_ net303 VGND VGND VPWR VPWR u_rf.reg31_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_38 _03282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 _01648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08170_ _03300_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__clkbuf_16
XANTENNA_27 _03176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07121_ _01606_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_49 _03320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_31_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_121_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_121_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_280 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput101 net101 VGND VGND VPWR VPWR adr_o[0] sky130_fd_sc_hd__buf_2
X_07052_ _01422_ _02251_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06003_ _01263_ _01266_ _01270_ _01273_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__nand4_1
Xoutput123 net123 VGND VGND VPWR VPWR adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput134 net134 VGND VGND VPWR VPWR icache_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput112 net112 VGND VGND VPWR VPWR adr_o[1] sky130_fd_sc_hd__buf_4
XFILLER_0_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput167 net167 VGND VGND VPWR VPWR store_data_o[0] sky130_fd_sc_hd__buf_4
Xoutput156 net156 VGND VGND VPWR VPWR icache_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput145 net145 VGND VGND VPWR VPWR icache_adr_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput178 net178 VGND VGND VPWR VPWR store_data_o[1] sky130_fd_sc_hd__clkbuf_4
Xoutput189 net189 VGND VGND VPWR VPWR store_data_o[2] sky130_fd_sc_hd__clkbuf_4
X_07954_ _03152_ _03161_ _02359_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_145_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07885_ _01272_ _01429_ _03095_ _01271_ VGND VGND VPWR VPWR _03096_ sky130_fd_sc_hd__o2bb2a_1
X_06905_ _02134_ _01437_ _02135_ _02155_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__a31oi_2
X_06836_ _02085_ _02089_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__nor2_2
X_09624_ u_rf.reg3_q\[16\] _04461_ _04582_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06767_ u_rf.reg0_q\[7\] _01516_ _01585_ u_rf.reg1_q\[7\] VGND VGND VPWR VPWR _02023_
+ sky130_fd_sc_hd__a22o_1
X_09555_ _04551_ VGND VGND VPWR VPWR _00080_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09486_ _04514_ VGND VGND VPWR VPWR _00048_ sky130_fd_sc_hd__clkbuf_1
X_08506_ u_rf.reg8_q\[16\] _03271_ _03273_ u_rf.reg29_q\[16\] _03693_ VGND VGND VPWR
+ VPWR _03694_ sky130_fd_sc_hd__a221o_1
X_06698_ _01450_ _01749_ _01956_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__a21o_1
X_08437_ u_rf.reg18_q\[13\] _03352_ _03348_ u_rf.reg9_q\[13\] _03627_ VGND VGND VPWR
+ VPWR _03628_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_186 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08368_ _03551_ _03562_ _03337_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__o21a_1
XFILLER_0_151_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08299_ _03480_ _03487_ _03496_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__or3_1
X_07319_ u_rf.reg3_q\[18\] _01606_ _01639_ u_rf.reg21_q\[18\] _02552_ VGND VGND VPWR
+ VPWR _02553_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_112_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_112_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10330_ u_rf.reg12_q\[27\] _04995_ _04981_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_429 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10261_ u_decod.rf_ff_res_data_i\[5\] VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__buf_2
X_12000_ clknet_leaf_83_clk u_exe.bu_pc_res\[13\] net365 VGND VGND VPWR VPWR u_exe.pc_data_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ _04738_ u_rf.reg11_q\[8\] _04900_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__mux2_1
Xfanout350 net351 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_2
Xfanout361 net367 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_4
XFILLER_0_17_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ clknet_leaf_140_clk _00939_ net204 VGND VGND VPWR VPWR u_rf.reg29_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12833_ clknet_leaf_118_clk _00870_ net326 VGND VGND VPWR VPWR u_rf.reg27_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12764_ clknet_leaf_127_clk _00801_ net238 VGND VGND VPWR VPWR u_rf.reg25_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11715_ clknet_leaf_129_clk _00007_ net234 VGND VGND VPWR VPWR u_rf.reg2_q\[7\] sky130_fd_sc_hd__dfrtp_1
X_12695_ clknet_leaf_70_clk _00732_ net352 VGND VGND VPWR VPWR u_rf.reg22_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_819 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11646_ u_decod.branch_imm_q_o\[2\] _01774_ _05696_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _04726_ u_rf.reg31_q\[2\] _05657_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__mux2_1
Xinput36 load_data_i[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput14 icache_instr_i[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
Xinput25 icache_instr_i[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_103_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_103_clk sky130_fd_sc_hd__clkbuf_16
X_10528_ _04768_ u_rf.reg15_q\[22\] _05100_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__mux2_1
Xinput69 reset_adr_i[13] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
Xinput58 load_data_i[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
Xinput47 load_data_i[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10459_ _05066_ VGND VGND VPWR VPWR _00469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12129_ clknet_leaf_117_clk _00166_ net326 VGND VGND VPWR VPWR u_rf.reg5_q\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07670_ u_rf.reg12_q\[25\] _01609_ _01628_ u_rf.reg29_q\[25\] _02889_ VGND VGND VPWR
+ VPWR _02890_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06621_ _01876_ _01878_ _01880_ _01882_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_36_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ _04409_ u_decod.rs2_data_q\[31\] _04410_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__and3_1
X_06552_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__or2_1
X_09271_ u_decod.pc_q_o\[31\] u_decod.branch_imm_q_o\[31\] VGND VGND VPWR VPWR _04382_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08222_ u_rf.reg0_q\[3\] _03420_ _03421_ u_rf.reg12_q\[3\] _03422_ VGND VGND VPWR
+ VPWR _03423_ sky130_fd_sc_hd__a221o_1
X_06483_ _01464_ _01749_ _01500_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08153_ _03264_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__buf_8
XFILLER_0_71_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07104_ _01950_ _02346_ _01467_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__mux2_1
X_08084_ u_rf.reg30_q\[0\] _03281_ _03283_ u_rf.reg10_q\[0\] _03287_ VGND VGND VPWR
+ VPWR _03288_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07035_ _02278_ _02280_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[12\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_58_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08986_ _04101_ _04136_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__nor2_1
X_07937_ u_rf.reg9_q\[31\] _02360_ _01668_ u_rf.reg8_q\[31\] _03144_ VGND VGND VPWR
+ VPWR _03145_ sky130_fd_sc_hd__a221o_1
X_07868_ u_decod.rf_ff_res_data_i\[29\] _02358_ _02743_ _03060_ _03079_ VGND VGND
+ VPWR VPWR _03080_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07799_ _02918_ _03013_ _01477_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
X_09607_ u_rf.reg3_q\[8\] _04444_ _04571_ VGND VGND VPWR VPWR _04580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06819_ u_rf.reg16_q\[8\] _01563_ _01629_ u_rf.reg17_q\[8\] VGND VGND VPWR VPWR _02073_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09538_ _04542_ VGND VGND VPWR VPWR _00072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_148_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ _05618_ VGND VGND VPWR VPWR _00958_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09469_ _04505_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_540 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ clknet_leaf_116_clk _00517_ net324 VGND VGND VPWR VPWR u_rf.reg16_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11431_ u_rf.reg28_q\[30\] u_decod.rf_ff_res_data_i\[30\] _05548_ VGND VGND VPWR
+ VPWR _05582_ sky130_fd_sc_hd__mux2_1
X_11362_ _05545_ VGND VGND VPWR VPWR _00893_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_78_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10313_ _04984_ VGND VGND VPWR VPWR _00405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11293_ u_rf.reg26_q\[29\] u_decod.rf_ff_res_data_i\[29\] _05499_ VGND VGND VPWR
+ VPWR _05509_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_60_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_91_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10244_ u_decod.rf_ff_rd_adr_q_i\[0\] _04424_ _04936_ VGND VGND VPWR VPWR _04937_
+ sky130_fd_sc_hd__or3_2
X_10175_ _04899_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12816_ clknet_leaf_34_clk _00853_ net275 VGND VGND VPWR VPWR u_rf.reg26_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_771 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12747_ clknet_leaf_135_clk _00784_ net208 VGND VGND VPWR VPWR u_rf.reg24_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12678_ clknet_leaf_140_clk _00715_ net204 VGND VGND VPWR VPWR u_rf.reg22_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11629_ _04778_ u_rf.reg31_q\[27\] _05679_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_100_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08840_ _03998_ _04011_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__nor2_1
XFILLER_0_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08771_ u_rf.reg1_q\[28\] _03310_ _03312_ u_rf.reg14_q\[28\] VGND VGND VPWR VPWR
+ _03947_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05983_ _01234_ _01074_ _01078_ _01252_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__and4_1
X_07722_ u_rf.reg16_q\[26\] _01565_ _02652_ u_rf.reg23_q\[26\] VGND VGND VPWR VPWR
+ _02940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_108_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07653_ u_decod.rs1_data_q\[25\] _01380_ u_decod.rs1_data_q\[9\] net377 _01468_ _01466_
+ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06604_ _01706_ _01750_ _01825_ _01866_ _01479_ _01476_ VGND VGND VPWR VPWR _01867_
+ sky130_fd_sc_hd__mux4_1
X_07584_ u_rf.reg1_q\[23\] _02604_ _01659_ u_rf.reg14_q\[23\] VGND VGND VPWR VPWR
+ _02808_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09323_ _01427_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_157_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06535_ _01779_ _01790_ _01800_ _01680_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09254_ u_decod.pc_q_o\[28\] u_decod.branch_imm_q_o\[28\] VGND VGND VPWR VPWR _04368_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06466_ u_rf.reg11_q\[1\] _01583_ _01638_ u_rf.reg21_q\[1\] _01733_ VGND VGND VPWR
+ VPWR _01734_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09185_ _04296_ _04303_ _04301_ _04300_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__a31o_1
X_08205_ net391 _03259_ _03406_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_554 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08136_ _03178_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__clkbuf_4
X_06397_ _01666_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_8
X_08067_ _03270_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07018_ u_rf.reg5_q\[12\] _01568_ _01555_ u_rf.reg6_q\[12\] VGND VGND VPWR VPWR _02264_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_126_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08969_ _04108_ _04111_ _04114_ _04121_ VGND VGND VPWR VPWR _04122_ sky130_fd_sc_hd__o31a_1
X_11980_ clknet_leaf_75_clk net451 net357 VGND VGND VPWR VPWR u_decod.pc_q_o\[29\]
+ sky130_fd_sc_hd__dfrtp_2
X_10931_ _05317_ VGND VGND VPWR VPWR _00690_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10862_ _05280_ VGND VGND VPWR VPWR _00658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12601_ clknet_leaf_62_clk _00638_ net343 VGND VGND VPWR VPWR u_rf.reg19_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10793_ u_rf.reg19_q\[18\] _04976_ _05235_ VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12532_ clknet_leaf_32_clk _00569_ net262 VGND VGND VPWR VPWR u_rf.reg17_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_774 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12463_ clknet_leaf_37_clk _00500_ net273 VGND VGND VPWR VPWR u_rf.reg15_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11414_ _05573_ VGND VGND VPWR VPWR _00917_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_671 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12394_ clknet_leaf_33_clk _00431_ net269 VGND VGND VPWR VPWR u_rf.reg13_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11345_ _04766_ u_rf.reg27_q\[21\] _05535_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11276_ _05500_ VGND VGND VPWR VPWR _00852_ sky130_fd_sc_hd__clkbuf_1
X_10227_ _04927_ VGND VGND VPWR VPWR _00376_ sky130_fd_sc_hd__clkbuf_1
X_13015_ clknet_leaf_66_clk _01052_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[28\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10158_ _04890_ VGND VGND VPWR VPWR _00344_ sky130_fd_sc_hd__clkbuf_1
X_10089_ u_rf.reg9_q\[24\] _04478_ _04849_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_832 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_638 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06320_ _01572_ _01515_ _01553_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__and3_2
XFILLER_0_155_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06251_ u_decod.exe_ff_rd_adr_q_i\[1\] VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06182_ u_decod.rs1_data_q\[5\] u_decod.rs1_data_q\[13\] _01358_ u_decod.rs1_data_q\[29\]
+ _01444_ _01447_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09941_ _04770_ u_rf.reg7_q\[23\] _04764_ VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap199 _02085_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_2
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ u_decod.rf_ff_res_data_i\[1\] VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__buf_2
X_08823_ u_decod.exe_ff_res_data_i\[30\] _03381_ _03996_ VGND VGND VPWR VPWR _03997_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08754_ u_rf.reg28_q\[27\] _03556_ _03557_ u_rf.reg2_q\[27\] VGND VGND VPWR VPWR
+ _03931_ sky130_fd_sc_hd__a22o_1
X_05966_ _01086_ _01087_ _01091_ VGND VGND VPWR VPWR _01244_ sky130_fd_sc_hd__and3_1
XFILLER_0_31_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07705_ _01481_ _02872_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08685_ u_rf.reg28_q\[24\] _03330_ _03332_ u_rf.reg2_q\[24\] VGND VGND VPWR VPWR
+ _03865_ sky130_fd_sc_hd__a22o_1
X_05897_ u_decod.pc0_q_i\[29\] _01186_ _01099_ VGND VGND VPWR VPWR _01190_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_92_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07636_ u_rf.reg5_q\[24\] _02664_ _01776_ u_rf.reg2_q\[24\] _02857_ VGND VGND VPWR
+ VPWR _02858_ sky130_fd_sc_hd__a221o_1
X_07567_ _02332_ _02771_ _02772_ _02791_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[23\]
+ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_24_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06518_ _01622_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__buf_6
XFILLER_0_91_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09306_ _04397_ u_decod.rs2_data_q\[15\] _04398_ VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09237_ _04345_ _04348_ _04346_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__a21boi_1
X_07498_ _01469_ _02346_ _01498_ VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_690 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06449_ u_decod.rf_ff_res_data_i\[1\] _01549_ _01714_ _01716_ VGND VGND VPWR VPWR
+ _01717_ sky130_fd_sc_hd__a22o_1
X_09168_ _04083_ _04274_ _04275_ _04294_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[15\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_90_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_384 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08119_ _03322_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__buf_6
XFILLER_0_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09099_ _04226_ u_decod.branch_imm_q_o\[4\] u_decod.pc_q_o\[4\] VGND VGND VPWR VPWR
+ _04235_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11130_ net527 _04972_ _05416_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11061_ _05386_ VGND VGND VPWR VPWR _00751_ sky130_fd_sc_hd__clkbuf_1
X_10012_ u_rf.reg8_q\[20\] _04469_ _04812_ VGND VGND VPWR VPWR _04813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
X_11963_ clknet_leaf_84_clk net459 net366 VGND VGND VPWR VPWR u_decod.pc_q_o\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11894_ clknet_leaf_96_clk u_decod.rs2_data_nxt\[15\] net333 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_10914_ u_rf.reg21_q\[10\] _04959_ _05308_ VGND VGND VPWR VPWR _05309_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_143_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10845_ u_rf.reg20_q\[10\] _04959_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10776_ _05223_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__buf_6
XFILLER_0_26_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12515_ clknet_leaf_110_clk _00552_ net315 VGND VGND VPWR VPWR u_rf.reg17_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12446_ clknet_leaf_136_clk _00483_ net205 VGND VGND VPWR VPWR u_rf.reg15_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12377_ clknet_leaf_58_clk _00414_ net292 VGND VGND VPWR VPWR u_rf.reg12_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11328_ _04749_ u_rf.reg27_q\[13\] _05524_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_152_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ _05491_ VGND VGND VPWR VPWR _00844_ sky130_fd_sc_hd__clkbuf_1
X_05820_ net468 _01105_ _01101_ net66 _01131_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__a221o_1
XFILLER_0_89_310 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
X_05751_ _01073_ VGND VGND VPWR VPWR _01074_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_148_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08470_ u_rf.reg27_q\[14\] _03318_ _03320_ u_rf.reg19_q\[14\] _03659_ VGND VGND VPWR
+ VPWR _03660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07421_ u_rf.reg12_q\[20\] _01609_ _01650_ u_rf.reg4_q\[20\] _02650_ VGND VGND VPWR
+ VPWR _02651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07352_ _02294_ _02400_ _02498_ _02584_ _01475_ _01905_ VGND VGND VPWR VPWR _02585_
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_359 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06303_ u_decod.dec0.instr_i\[22\] _01537_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__nor2_2
XFILLER_0_116_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07283_ u_rf.reg3_q\[17\] _01605_ _01638_ u_rf.reg21_q\[17\] _02518_ VGND VGND VPWR
+ VPWR _02519_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_150_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_805 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09022_ u_decod.rs1_data_q\[30\] u_decod.branch_imm_q_o\[30\] VGND VGND VPWR VPWR
+ _04167_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06234_ _01504_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06165_ u_decod.instr_unit_q\[0\] u_decod.instr_operation_q\[0\] _01427_ VGND VGND
+ VPWR VPWR _01436_ sky130_fd_sc_hd__and3_2
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06096_ u_decod.rs1_data_q\[23\] VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09924_ u_decod.rf_ff_res_data_i\[18\] VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09855_ _04713_ VGND VGND VPWR VPWR _00218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08806_ u_rf.reg31_q\[30\] _03289_ _03291_ u_rf.reg11_q\[30\] _03979_ VGND VGND VPWR
+ VPWR _03980_ sky130_fd_sc_hd__a221o_1
X_09786_ _04676_ VGND VGND VPWR VPWR _00186_ sky130_fd_sc_hd__clkbuf_1
X_06998_ _01763_ _02244_ _01298_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ u_decod.exe_ff_res_data_i\[26\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[26\]
+ _03914_ VGND VGND VPWR VPWR _03915_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_65_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_106 u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05949_ _01227_ _01229_ VGND VGND VPWR VPWR _01230_ sky130_fd_sc_hd__or2_1
X_08668_ u_rf.reg16_q\[23\] _03450_ _03515_ u_rf.reg5_q\[23\] VGND VGND VPWR VPWR
+ _03849_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 _01605_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_117 u_rf.reg8_q\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 _02002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ _01572_ _01224_ _02646_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__a21o_2
X_08599_ u_rf.reg6_q\[20\] _03305_ _03307_ u_rf.reg13_q\[20\] VGND VGND VPWR VPWR
+ _03783_ sky130_fd_sc_hd__a22o_1
X_10630_ u_rf.reg17_q\[5\] _04949_ _05152_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_284 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10561_ _05121_ VGND VGND VPWR VPWR _00516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_608 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12300_ clknet_leaf_9_clk _00337_ net266 VGND VGND VPWR VPWR u_rf.reg10_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_10492_ _04732_ u_rf.reg15_q\[5\] _05078_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12231_ clknet_leaf_4_clk _00268_ net211 VGND VGND VPWR VPWR u_rf.reg8_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12162_ clknet_leaf_131_clk _00199_ net229 VGND VGND VPWR VPWR u_rf.reg6_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12093_ clknet_leaf_15_clk _00130_ net245 VGND VGND VPWR VPWR u_rf.reg4_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_11113_ u_rf.reg24_q\[8\] _04955_ _05405_ VGND VGND VPWR VPWR _05414_ sky130_fd_sc_hd__mux2_1
X_11044_ _05377_ VGND VGND VPWR VPWR _00743_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ clknet_leaf_92_clk _01032_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[8\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11946_ clknet_leaf_115_clk u_decod.dec0.rd_o\[0\] net328 VGND VGND VPWR VPWR u_decod.exe_ff_rd_adr_q_i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11877_ clknet_leaf_103_clk u_decod.dec0.access_size_o\[1\] net335 VGND VGND VPWR
+ VPWR net99 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10828_ u_rf.reg20_q\[2\] _04943_ _05260_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10759_ _05226_ VGND VGND VPWR VPWR _00609_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_12 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12429_ clknet_leaf_5_clk _00466_ net217 VGND VGND VPWR VPWR u_rf.reg14_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_381 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07970_ _03175_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__buf_6
XFILLER_0_10_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06921_ u_rf.reg13_q\[10\] _01596_ _01590_ u_rf.reg18_q\[10\] _02170_ VGND VGND VPWR
+ VPWR _02171_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_147_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_147_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09640_ _04597_ VGND VGND VPWR VPWR _00119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06852_ net64 _02047_ _02049_ net50 _02051_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__a221oi_1
X_05803_ _01100_ VGND VGND VPWR VPWR _01119_ sky130_fd_sc_hd__clkbuf_4
X_09571_ u_rf.reg0_q\[24\] _04478_ _04555_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__mux2_1
X_06783_ u_decod.rs1_data_q\[23\] _01683_ u_decod.rs1_data_q\[15\] _01267_ _01445_
+ _01684_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_47_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_05734_ u_decod.branch_imm_q_o\[1\] u_decod.rs1_data_q\[1\] VGND VGND VPWR VPWR _01060_
+ sky130_fd_sc_hd__xor2_2
XFILLER_0_78_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08522_ u_decod.exe_ff_res_data_i\[16\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[16\]
+ _03709_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08453_ _03637_ _03639_ _03641_ _03643_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__or4_1
XFILLER_0_78_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07404_ _02411_ _01293_ _02331_ _01392_ _01291_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__a311o_1
XFILLER_0_147_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08384_ u_rf.reg7_q\[10\] _03428_ _03429_ u_rf.reg25_q\[10\] _03577_ VGND VGND VPWR
+ VPWR _03578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07335_ _02562_ _02564_ _02566_ _02568_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_63_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07266_ _01383_ _02244_ _01431_ _01382_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09005_ _04132_ _04139_ _04144_ _04149_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06217_ net112 _01066_ _01486_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__and3_2
XFILLER_0_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07197_ _02430_ _02432_ _02434_ _02436_ VGND VGND VPWR VPWR _02437_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06148_ u_decod.rs2_data_q\[32\] u_decod.rs1_data_q\[32\] VGND VGND VPWR VPWR _01419_
+ sky130_fd_sc_hd__xnor2_4
X_06079_ _01348_ _01349_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__nor2_1
X_09907_ _04747_ u_rf.reg7_q\[12\] _04743_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__mux2_1
X_09838_ _04704_ VGND VGND VPWR VPWR _00210_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09769_ _04667_ VGND VGND VPWR VPWR _00178_ sky130_fd_sc_hd__clkbuf_1
X_11800_ clknet_leaf_76_clk net153 net369 VGND VGND VPWR VPWR u_decod.pc0_q_i\[27\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_38_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_83_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12780_ clknet_leaf_20_clk _00817_ net280 VGND VGND VPWR VPWR u_rf.reg25_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_83_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11731_ clknet_leaf_41_clk _00023_ net277 VGND VGND VPWR VPWR u_rf.reg2_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11662_ net518 _05700_ _02644_ _05705_ VGND VGND VPWR VPWR _01033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10613_ _05148_ VGND VGND VPWR VPWR _00541_ sky130_fd_sc_hd__clkbuf_1
X_11593_ _05656_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_12_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_221 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10544_ _04784_ u_rf.reg15_q\[30\] _05077_ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10475_ _05074_ VGND VGND VPWR VPWR _00477_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_114_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12214_ clknet_leaf_48_clk _00251_ net306 VGND VGND VPWR VPWR u_rf.reg7_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_156 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12145_ clknet_leaf_55_clk _00182_ net284 VGND VGND VPWR VPWR u_rf.reg5_q\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12076_ clknet_leaf_26_clk _00113_ net266 VGND VGND VPWR VPWR u_rf.reg3_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_11027_ _01532_ _01536_ _04568_ _05114_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__or4_4
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
X_12978_ clknet_leaf_46_clk _01015_ net299 VGND VGND VPWR VPWR u_rf.reg31_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11929_ clknet_leaf_101_clk u_decod.rs1_data\[17\] net338 VGND VGND VPWR VPWR u_decod.rs1_data_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_210 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _01650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_28 _03200_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_39 _03283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07120_ u_rf.reg0_q\[14\] _01664_ _02360_ u_rf.reg9_q\[14\] _02361_ VGND VGND VPWR
+ VPWR _02362_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07051_ _02292_ _02295_ _01474_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput113 net113 VGND VGND VPWR VPWR adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput124 net124 VGND VGND VPWR VPWR adr_o[30] sky130_fd_sc_hd__buf_6
XFILLER_0_112_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06002_ _01271_ _01272_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput102 net102 VGND VGND VPWR VPWR adr_o[10] sky130_fd_sc_hd__buf_2
XFILLER_0_3_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput146 net146 VGND VGND VPWR VPWR icache_adr_o[20] sky130_fd_sc_hd__buf_2
Xoutput157 net157 VGND VGND VPWR VPWR icache_adr_o[30] sky130_fd_sc_hd__buf_6
Xoutput135 net135 VGND VGND VPWR VPWR icache_adr_o[10] sky130_fd_sc_hd__buf_4
XFILLER_0_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput168 net168 VGND VGND VPWR VPWR store_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput179 net179 VGND VGND VPWR VPWR store_data_o[20] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_699 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07953_ _03154_ _03156_ _03158_ _03160_ VGND VGND VPWR VPWR _03161_ sky130_fd_sc_hd__or4_1
X_07884_ _01272_ _02244_ _01820_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__o21a_1
X_06904_ _01441_ _02140_ _02147_ _02154_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09623_ _04588_ VGND VGND VPWR VPWR _00111_ sky130_fd_sc_hd__clkbuf_1
X_06835_ _02088_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_39_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06766_ _02015_ _02017_ _02019_ _02021_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__or4_1
X_09554_ u_rf.reg0_q\[16\] _04461_ _04544_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09485_ u_rf.reg1_q\[16\] _04461_ _04507_ VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__mux2_1
X_08505_ u_rf.reg22_q\[16\] _03409_ _03277_ u_rf.reg3_q\[16\] VGND VGND VPWR VPWR
+ _03693_ sky130_fd_sc_hd__a22o_1
X_06697_ u_decod.rs2_data_q\[3\] _01955_ _01497_ _01457_ VGND VGND VPWR VPWR _01956_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08436_ u_rf.reg29_q\[13\] _03217_ _03213_ u_rf.reg20_q\[13\] VGND VGND VPWR VPWR
+ _03627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_850 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08367_ _03553_ _03555_ _03559_ _03561_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__or4_1
XFILLER_0_74_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07318_ u_rf.reg5_q\[18\] _01568_ _01556_ u_rf.reg6_q\[18\] VGND VGND VPWR VPWR _02552_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08298_ _03489_ _03491_ _03493_ _03495_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__or4_1
XFILLER_0_144_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07249_ _02394_ _02395_ _02440_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__and3b_2
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10260_ _04948_ VGND VGND VPWR VPWR _00388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10191_ _04908_ VGND VGND VPWR VPWR _00359_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_874 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout340 net348 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_4
Xfanout351 net359 VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_4
Xfanout373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_4
Xfanout362 net367 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_4
X_12901_ clknet_leaf_125_clk _00938_ net240 VGND VGND VPWR VPWR u_rf.reg29_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12832_ clknet_leaf_120_clk _00869_ net249 VGND VGND VPWR VPWR u_rf.reg27_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ clknet_leaf_13_clk _00800_ net244 VGND VGND VPWR VPWR u_rf.reg25_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11714_ clknet_leaf_16_clk _00006_ net250 VGND VGND VPWR VPWR u_rf.reg2_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_316 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12694_ clknet_leaf_49_clk _00731_ net307 VGND VGND VPWR VPWR u_rf.reg22_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_749 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11645_ net355 VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput37 load_data_i[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
XFILLER_0_52_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput15 icache_instr_i[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
Xinput26 icache_instr_i[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
X_11576_ _05659_ VGND VGND VPWR VPWR _00993_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10527_ _05102_ VGND VGND VPWR VPWR _00501_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput59 load_data_i[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
Xinput48 load_data_i[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10458_ _04766_ u_rf.reg14_q\[21\] _05064_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10389_ _05029_ VGND VGND VPWR VPWR _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12128_ clknet_leaf_121_clk _00165_ net247 VGND VGND VPWR VPWR u_rf.reg5_q\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12059_ clknet_leaf_11_clk _00096_ net221 VGND VGND VPWR VPWR u_rf.reg3_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_06620_ u_rf.reg29_q\[4\] _01628_ _01638_ u_rf.reg21_q\[4\] _01881_ VGND VGND VPWR
+ VPWR _01882_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_140_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_36_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06551_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_47_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_305 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09270_ _04197_ _04380_ _04381_ _04200_ _04170_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[30\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_114_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06482_ _01444_ _01748_ _01497_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08221_ u_rf.reg28_q\[3\] _03330_ _03332_ u_rf.reg2_q\[3\] VGND VGND VPWR VPWR _03422_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08152_ _03354_ VGND VGND VPWR VPWR _03355_ sky130_fd_sc_hd__buf_8
XFILLER_0_16_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07103_ u_decod.rs1_data_q\[29\] _01447_ _02136_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__o21a_1
X_08083_ u_rf.reg26_q\[0\] _03284_ _03286_ u_rf.reg21_q\[0\] VGND VGND VPWR VPWR _03287_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07034_ _01897_ _02279_ _02090_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08985_ _04132_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07936_ u_rf.reg30_q\[31\] _01581_ _02419_ u_rf.reg28_q\[31\] VGND VGND VPWR VPWR
+ _03144_ sky130_fd_sc_hd__a22o_1
X_07867_ _03069_ _03078_ _02359_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__o21a_1
XFILLER_0_155_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07798_ _02833_ _03012_ _02685_ VGND VGND VPWR VPWR _03013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09606_ _04579_ VGND VGND VPWR VPWR _00103_ sky130_fd_sc_hd__clkbuf_1
X_06818_ _02065_ _02067_ _02069_ _02071_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09537_ u_rf.reg0_q\[8\] _04444_ _04533_ VGND VGND VPWR VPWR _04542_ sky130_fd_sc_hd__mux2_1
X_06749_ u_decod.pc_q_o\[6\] u_decod.pc_q_o\[7\] _01917_ VGND VGND VPWR VPWR _02006_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_65_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09468_ u_rf.reg1_q\[8\] _04444_ _04496_ VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09399_ _04460_ VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__clkbuf_1
X_08419_ u_rf.reg9_q\[12\] _03348_ _03349_ u_rf.reg20_q\[12\] VGND VGND VPWR VPWR
+ _03611_ sky130_fd_sc_hd__a22o_1
X_11430_ _05581_ VGND VGND VPWR VPWR _00925_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11361_ _04782_ u_rf.reg27_q\[29\] _05535_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_363 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10312_ u_rf.reg12_q\[21\] _04983_ _04981_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11292_ _05508_ VGND VGND VPWR VPWR _00860_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10243_ _01531_ _01536_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__nand2_2
X_10174_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12815_ clknet_leaf_42_clk _00852_ net276 VGND VGND VPWR VPWR u_rf.reg26_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_351 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12746_ clknet_leaf_30_clk _00783_ net261 VGND VGND VPWR VPWR u_rf.reg24_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12677_ clknet_leaf_125_clk _00714_ net239 VGND VGND VPWR VPWR u_rf.reg22_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11628_ _05686_ VGND VGND VPWR VPWR _01018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11559_ _04776_ u_rf.reg30_q\[26\] _05643_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08770_ u_rf.reg15_q\[28\] _03373_ _03374_ u_rf.reg24_q\[28\] _03945_ VGND VGND VPWR
+ VPWR _03946_ sky130_fd_sc_hd__a221o_1
X_05982_ _01255_ VGND VGND VPWR VPWR u_decod.dec0.access_size_o\[1\] sky130_fd_sc_hd__clkbuf_1
X_07721_ _02932_ _02934_ _02936_ _02938_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07652_ _02830_ _02872_ _01425_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07583_ u_rf.reg25_q\[23\] _01783_ _01784_ u_rf.reg24_q\[23\] _02806_ VGND VGND VPWR
+ VPWR _02807_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06603_ _01499_ _01865_ _01458_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09322_ u_decod.instr_unit_q\[3\] VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__buf_2
X_06534_ _01793_ _01795_ _01797_ _01799_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09253_ _04362_ _04365_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__nand3_1
XFILLER_0_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06465_ u_rf.reg15_q\[1\] _01600_ _01608_ u_rf.reg12_q\[1\] VGND VGND VPWR VPWR _01733_
+ sky130_fd_sc_hd__a22o_1
X_09184_ _04306_ _04307_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__nand2_1
X_08204_ u_decod.exe_ff_res_data_i\[2\] _03381_ _03405_ VGND VGND VPWR VPWR _03406_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_62_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06396_ _01665_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08135_ u_decod.exe_ff_res_data_i\[0\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[0\]
+ _03338_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08066_ _03216_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__clkbuf_8
X_07017_ u_rf.reg0_q\[12\] _01663_ _01636_ u_rf.reg9_q\[12\] _02262_ VGND VGND VPWR
+ VPWR _02263_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_73_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08968_ _01358_ u_decod.branch_imm_q_o\[21\] _04120_ VGND VGND VPWR VPWR _04121_
+ sky130_fd_sc_hd__a21oi_1
X_08899_ _04060_ _04061_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__nor2_1
X_07919_ _01273_ _03083_ _01272_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a21oi_1
X_10930_ u_rf.reg21_q\[18\] _04976_ _05308_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__mux2_1
X_12600_ clknet_leaf_63_clk _00637_ net342 VGND VGND VPWR VPWR u_rf.reg19_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10861_ u_rf.reg20_q\[18\] _04976_ _05271_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10792_ _05243_ VGND VGND VPWR VPWR _00625_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_455 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12531_ clknet_leaf_53_clk _00568_ net305 VGND VGND VPWR VPWR u_rf.reg17_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12462_ clknet_leaf_27_clk _00499_ net258 VGND VGND VPWR VPWR u_rf.reg15_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11413_ u_rf.reg28_q\[21\] u_decod.rf_ff_res_data_i\[21\] _05571_ VGND VGND VPWR
+ VPWR _05573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12393_ clknet_leaf_56_clk _00430_ net286 VGND VGND VPWR VPWR u_rf.reg13_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_571 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11344_ _05536_ VGND VGND VPWR VPWR _00884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11275_ u_rf.reg26_q\[20\] u_decod.rf_ff_res_data_i\[20\] _05499_ VGND VGND VPWR
+ VPWR _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13014_ clknet_leaf_74_clk _01051_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[27\]
+ sky130_fd_sc_hd__dfxtp_1
X_10226_ _04772_ u_rf.reg11_q\[24\] _04922_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__mux2_1
X_10157_ u_rf.reg10_q\[24\] _04478_ _04885_ VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10088_ _04853_ VGND VGND VPWR VPWR _00311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12729_ clknet_leaf_63_clk _00766_ net342 VGND VGND VPWR VPWR u_rf.reg23_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06250_ u_decod.dec0.instr_i\[20\] VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__inv_2
XFILLER_0_155_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06181_ _01448_ _01449_ _01451_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09940_ u_decod.rf_ff_res_data_i\[23\] VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__buf_2
XFILLER_0_111_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09871_ _04723_ VGND VGND VPWR VPWR _00224_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ u_decod.rf_ff_res_data_i\[30\] _03197_ _03995_ _03404_ VGND VGND VPWR VPWR
+ _03996_ sky130_fd_sc_hd__a22o_1
X_08753_ u_rf.reg27_q\[27\] _03365_ _03366_ u_rf.reg19_q\[27\] _03929_ VGND VGND VPWR
+ VPWR _03930_ sky130_fd_sc_hd__a221o_1
X_05965_ u_decod.dec0.funct3\[2\] _01241_ VGND VGND VPWR VPWR _01243_ sky130_fd_sc_hd__and2_2
X_07704_ _01481_ _02922_ _01443_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08684_ _03857_ _03859_ _03861_ _03863_ VGND VGND VPWR VPWR _03864_ sky130_fd_sc_hd__or4_1
X_05896_ u_decod.pc0_q_i\[29\] _01186_ VGND VGND VPWR VPWR _01189_ sky130_fd_sc_hd__and2_1
X_07635_ u_rf.reg15_q\[24\] _02371_ _02652_ u_rf.reg23_q\[24\] VGND VGND VPWR VPWR
+ _02857_ sky130_fd_sc_hd__a22o_1
X_07566_ _02775_ _02777_ _02784_ _02790_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__or4b_1
X_06517_ _01576_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__buf_6
X_09305_ _04400_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09236_ _04350_ _04351_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__nand2_1
X_07497_ _02624_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06448_ u_decod.dec0.instr_i\[8\] _01226_ _01715_ u_decod.dec0.instr_i\[21\] VGND
+ VGND VPWR VPWR _01716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09167_ _04292_ _04293_ VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__xnor2_1
X_06379_ _01648_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08118_ _03248_ VGND VGND VPWR VPWR _03322_ sky130_fd_sc_hd__buf_8
X_09098_ _04227_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08049_ u_decod.exe_ff_res_data_i\[31\] _03187_ _03197_ u_decod.rf_ff_res_data_i\[31\]
+ _03254_ VGND VGND VPWR VPWR _03255_ sky130_fd_sc_hd__a221o_1
X_11060_ _04753_ u_rf.reg23_q\[15\] _05380_ VGND VGND VPWR VPWR _05386_ sky130_fd_sc_hd__mux2_1
X_10011_ _04789_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11962_ clknet_leaf_85_clk net448 net362 VGND VGND VPWR VPWR u_decod.pc_q_o\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_86_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10913_ _05296_ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__buf_6
X_11893_ clknet_leaf_96_clk u_decod.rs2_data_nxt\[14\] net332 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10844_ _05259_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__buf_8
XFILLER_0_67_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12514_ clknet_leaf_133_clk _00551_ net231 VGND VGND VPWR VPWR u_rf.reg17_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10775_ _05234_ VGND VGND VPWR VPWR _00617_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_162 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_789 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12445_ clknet_leaf_15_clk _00482_ net245 VGND VGND VPWR VPWR u_rf.reg15_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_117_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12376_ clknet_leaf_63_clk _00413_ net342 VGND VGND VPWR VPWR u_rf.reg12_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11327_ _05527_ VGND VGND VPWR VPWR _00876_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11258_ u_rf.reg26_q\[12\] u_decod.rf_ff_res_data_i\[12\] _05488_ VGND VGND VPWR
+ VPWR _05491_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10209_ _04755_ u_rf.reg11_q\[16\] _04911_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__mux2_1
X_11189_ _05454_ VGND VGND VPWR VPWR _00811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05750_ u_decod.dec0.instr_i\[2\] u_decod.dec0.instr_i\[1\] _01072_ VGND VGND VPWR
+ VPWR _01073_ sky130_fd_sc_hd__and3b_1
XFILLER_0_82_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07420_ u_rf.reg31_q\[20\] _01616_ _01791_ u_rf.reg10_q\[20\] VGND VGND VPWR VPWR
+ _02650_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07351_ _01376_ u_decod.rs1_data_q\[11\] u_decod.rs1_data_q\[3\] _01747_ _01467_
+ _01461_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__mux4_2
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06302_ _01538_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_116_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07282_ u_rf.reg5_q\[17\] _01568_ _01555_ u_rf.reg6_q\[17\] VGND VGND VPWR VPWR _02518_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09021_ u_decod.rs1_data_q\[30\] u_decod.branch_imm_q_o\[30\] VGND VGND VPWR VPWR
+ _04166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06233_ u_decod.instr_operation_q\[0\] u_decod.instr_unit_q\[1\] _01427_ VGND VGND
+ VPWR VPWR _01504_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06164_ _01434_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__buf_4
XFILLER_0_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06095_ _01364_ _01365_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09923_ _04758_ VGND VGND VPWR VPWR _00241_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09854_ u_rf.reg6_q\[26\] _04482_ _04706_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08805_ u_rf.reg9_q\[30\] _03293_ _03295_ u_rf.reg20_q\[30\] VGND VGND VPWR VPWR
+ _03979_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09785_ u_rf.reg5_q\[26\] _04482_ _04669_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__mux2_1
X_06997_ _01697_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_29_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08736_ _03904_ _03913_ _03378_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__o21a_1
XANTENNA_107 u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_05948_ _01094_ _01228_ _01074_ _01092_ VGND VGND VPWR VPWR _01229_ sky130_fd_sc_hd__o211a_1
X_08667_ u_rf.reg7_q\[23\] _03428_ _03429_ u_rf.reg25_q\[23\] _03847_ VGND VGND VPWR
+ VPWR _03848_ sky130_fd_sc_hd__a221o_1
X_05879_ _01099_ _01174_ _01175_ _01176_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__a31o_1
XFILLER_0_96_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 _01610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_07618_ _02840_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[24\] sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_101_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08598_ _03775_ _03777_ _03779_ _03781_ VGND VGND VPWR VPWR _03782_ sky130_fd_sc_hd__or4_1
XFILLER_0_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07549_ u_decod.pc_q_o\[21\] u_decod.pc_q_o\[22\] _02638_ u_decod.pc_q_o\[23\] VGND
+ VGND VPWR VPWR _02774_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_81_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10560_ u_rf.reg16_q\[4\] _04947_ _05116_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09219_ _04328_ _04331_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10491_ _05083_ VGND VGND VPWR VPWR _00484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12230_ clknet_leaf_140_clk _00267_ net202 VGND VGND VPWR VPWR u_rf.reg8_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12161_ clknet_leaf_120_clk _00198_ net326 VGND VGND VPWR VPWR u_rf.reg6_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12092_ clknet_leaf_128_clk _00129_ net234 VGND VGND VPWR VPWR u_rf.reg4_q\[1\] sky130_fd_sc_hd__dfrtp_1
X_11112_ _05413_ VGND VGND VPWR VPWR _00775_ sky130_fd_sc_hd__clkbuf_1
X_11043_ _04736_ u_rf.reg23_q\[7\] _05369_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
X_12994_ clknet_leaf_92_clk _01031_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[7\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_87_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11945_ clknet_leaf_97_clk u_decod.dec0.rd_v net332 VGND VGND VPWR VPWR u_decod.rd_v_q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_539 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11876_ clknet_leaf_103_clk u_decod.dec0.access_size_o\[0\] net335 VGND VGND VPWR
+ VPWR net98 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_380 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10827_ _05262_ VGND VGND VPWR VPWR _00641_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10758_ u_rf.reg19_q\[1\] _04941_ _05224_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12428_ clknet_leaf_19_clk _00465_ net281 VGND VGND VPWR VPWR u_rf.reg14_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ _05189_ VGND VGND VPWR VPWR _00576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12359_ clknet_leaf_4_clk _00396_ net212 VGND VGND VPWR VPWR u_rf.reg12_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06920_ u_rf.reg30_q\[10\] _01578_ _01623_ u_rf.reg28_q\[10\] VGND VGND VPWR VPWR
+ _02170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_147_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06851_ _01478_ _02102_ _02103_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__o21ai_1
X_09570_ _04559_ VGND VGND VPWR VPWR _00087_ sky130_fd_sc_hd__clkbuf_1
X_05802_ _01104_ VGND VGND VPWR VPWR _01118_ sky130_fd_sc_hd__buf_4
X_06782_ _02035_ _02037_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05733_ _01059_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_4
X_08521_ _03699_ _03708_ _03378_ VGND VGND VPWR VPWR _03709_ sky130_fd_sc_hd__o21a_2
XFILLER_0_148_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08452_ u_rf.reg30_q\[13\] _03280_ _03325_ u_rf.reg5_q\[13\] _03642_ VGND VGND VPWR
+ VPWR _03643_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07403_ _01442_ _02626_ _02628_ _02633_ VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_594 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08383_ u_rf.reg1_q\[10\] _03446_ _03447_ u_rf.reg14_q\[10\] VGND VGND VPWR VPWR
+ _03577_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07334_ u_rf.reg16_q\[18\] _01565_ _01674_ u_rf.reg2_q\[18\] _02567_ VGND VGND VPWR
+ VPWR _02568_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_63_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07265_ _01422_ _02499_ _02501_ _01505_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09004_ _04101_ _04151_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__nor2_1
XFILLER_0_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06216_ _01064_ _01067_ _01486_ net100 VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__a31o_2
X_07196_ u_rf.reg20_q\[15\] _02385_ _02386_ u_rf.reg27_q\[15\] _02435_ VGND VGND VPWR
+ VPWR _02436_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06147_ _01274_ _01413_ _01417_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__o21a_1
X_06078_ u_decod.rs2_data_q\[12\] _01297_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09906_ u_decod.rf_ff_res_data_i\[12\] VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09837_ u_rf.reg6_q\[18\] _04465_ _04695_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__mux2_1
X_09768_ u_rf.reg5_q\[18\] _04465_ _04658_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__mux2_1
X_08719_ u_rf.reg4_q\[26\] _03356_ _03357_ u_rf.reg17_q\[26\] _03896_ VGND VGND VPWR
+ VPWR _03897_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11730_ clknet_leaf_55_clk _00022_ net286 VGND VGND VPWR VPWR u_rf.reg2_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ u_rf.reg4_q\[19\] _04467_ _04619_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11661_ _05693_ u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10612_ net529 _04999_ _05138_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11592_ _05667_ VGND VGND VPWR VPWR _01001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_233 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10543_ _05110_ VGND VGND VPWR VPWR _00509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10474_ _04782_ u_rf.reg14_q\[29\] _05064_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12213_ clknet_leaf_47_clk _00250_ net300 VGND VGND VPWR VPWR u_rf.reg7_q\[26\] sky130_fd_sc_hd__dfrtp_1
X_12144_ clknet_leaf_32_clk _00181_ net263 VGND VGND VPWR VPWR u_rf.reg5_q\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_94_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12075_ clknet_leaf_1_clk _00112_ net208 VGND VGND VPWR VPWR u_rf.reg3_q\[16\] sky130_fd_sc_hd__dfrtp_1
X_11026_ _05367_ VGND VGND VPWR VPWR _00735_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ clknet_leaf_55_clk _01014_ net294 VGND VGND VPWR VPWR u_rf.reg31_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11928_ clknet_leaf_101_clk u_decod.rs1_data\[16\] net338 VGND VGND VPWR VPWR u_decod.rs1_data_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11859_ clknet_leaf_55_clk _00086_ net284 VGND VGND VPWR VPWR u_rf.reg0_q\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _01652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _03202_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_383 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07050_ _02094_ _02294_ _01458_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06001_ u_decod.rs2_data_q\[30\] u_decod.rs1_data_q\[30\] VGND VGND VPWR VPWR _01272_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_88_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR adr_o[21] sky130_fd_sc_hd__buf_4
Xoutput125 net125 VGND VGND VPWR VPWR adr_o[31] sky130_fd_sc_hd__buf_8
Xoutput103 net103 VGND VGND VPWR VPWR adr_o[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput147 net147 VGND VGND VPWR VPWR icache_adr_o[21] sky130_fd_sc_hd__buf_4
Xoutput158 net158 VGND VGND VPWR VPWR icache_adr_o[31] sky130_fd_sc_hd__clkbuf_4
Xoutput136 net136 VGND VGND VPWR VPWR icache_adr_o[11] sky130_fd_sc_hd__buf_6
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput169 net169 VGND VGND VPWR VPWR store_data_o[11] sky130_fd_sc_hd__clkbuf_4
X_07952_ u_rf.reg5_q\[31\] _02664_ _02665_ u_rf.reg19_q\[31\] _03159_ VGND VGND VPWR
+ VPWR _03160_ sky130_fd_sc_hd__a221o_1
X_07883_ _03089_ _03093_ _01481_ VGND VGND VPWR VPWR _03094_ sky130_fd_sc_hd__mux2_1
X_06903_ _01058_ _02148_ _02153_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__a21bo_1
X_09622_ u_rf.reg3_q\[15\] _04459_ _04582_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__mux2_1
X_06834_ _01804_ _02086_ _01898_ _02087_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__and4_1
X_09553_ _04550_ VGND VGND VPWR VPWR _00079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ u_rf.reg18_q\[16\] _03262_ _03263_ u_rf.reg23_q\[16\] _03691_ VGND VGND VPWR
+ VPWR _03692_ sky130_fd_sc_hd__a221o_1
X_06765_ u_rf.reg30_q\[7\] _01579_ _01655_ u_rf.reg10_q\[7\] _02020_ VGND VGND VPWR
+ VPWR _02021_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09484_ _04513_ VGND VGND VPWR VPWR _00047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06696_ u_decod.rs1_data_q\[6\] _01445_ _01703_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__o21a_1
X_08435_ u_decod.pc0_q_i\[12\] _03565_ _03626_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[12\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08366_ u_rf.reg16_q\[9\] _03323_ _03325_ u_rf.reg5_q\[9\] _03560_ VGND VGND VPWR
+ VPWR _03561_ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07317_ u_decod.dec0.instr_i\[18\] _01208_ _02256_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08297_ u_rf.reg18_q\[6\] _03352_ _03354_ u_rf.reg23_q\[6\] _03494_ VGND VGND VPWR
+ VPWR _03495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07248_ _01713_ u_decod.exe_ff_res_data_i\[16\] _02485_ VGND VGND VPWR VPWR _02486_
+ sky130_fd_sc_hd__a21o_1
X_07179_ _01625_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10190_ _04736_ u_rf.reg11_q\[7\] _04900_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout341 net348 VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_4
Xfanout330 net334 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__buf_2
Xfanout352 net354 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_4
Xfanout363 net367 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
Xfanout374 net97 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_8
X_12900_ clknet_leaf_107_clk _00937_ net315 VGND VGND VPWR VPWR u_rf.reg29_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12831_ clknet_leaf_137_clk _00868_ net206 VGND VGND VPWR VPWR u_rf.reg27_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ clknet_leaf_60_clk _00799_ net290 VGND VGND VPWR VPWR u_rf.reg24_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12693_ clknet_leaf_47_clk _00730_ net301 VGND VGND VPWR VPWR u_rf.reg22_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11713_ clknet_leaf_122_clk _00005_ net247 VGND VGND VPWR VPWR u_rf.reg2_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11644_ _05695_ VGND VGND VPWR VPWR _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 icache_instr_i[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 icache_instr_i[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
X_11575_ _04724_ u_rf.reg31_q\[1\] _05657_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10526_ _04766_ u_rf.reg15_q\[21\] _05100_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput49 load_data_i[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 load_data_i[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s2s_1
X_10457_ _05065_ VGND VGND VPWR VPWR _00468_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10388_ _04763_ u_rf.reg13_q\[20\] _05028_ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12127_ clknet_leaf_137_clk _00164_ net206 VGND VGND VPWR VPWR u_rf.reg5_q\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12058_ clknet_leaf_88_clk u_exe.branch_v net361 VGND VGND VPWR VPWR u_decod.flush_v
+ sky130_fd_sc_hd__dfrtp_4
X_11009_ u_rf.reg22_q\[23\] _04987_ _05355_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06550_ _01811_ _01813_ _01814_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_114 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06481_ _01445_ u_decod.rs1_data_q\[2\] _01703_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08220_ _03328_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__buf_6
XFILLER_0_145_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08151_ _03223_ VGND VGND VPWR VPWR _03354_ sky130_fd_sc_hd__buf_8
XFILLER_0_99_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08082_ _03285_ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__buf_8
X_07102_ _02239_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07033_ _02225_ _02226_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08984_ _04119_ _04122_ _04126_ _04134_ VGND VGND VPWR VPWR _04135_ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07935_ _01224_ _02644_ u_decod.dec0.funct7\[6\] VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_707 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07866_ _03071_ _03073_ _03075_ _03077_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09605_ u_rf.reg3_q\[7\] _04442_ _04571_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07797_ u_decod.rs1_data_q\[28\] _01363_ _01297_ u_decod.rs1_data_q\[4\] _01469_
+ _01466_ VGND VGND VPWR VPWR _03012_ sky130_fd_sc_hd__mux4_1
X_06817_ u_rf.reg12_q\[8\] _01607_ _01672_ u_rf.reg2_q\[8\] _02070_ VGND VGND VPWR
+ VPWR _02071_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06748_ u_decod.pc_q_o\[6\] _01917_ u_decod.pc_q_o\[7\] VGND VGND VPWR VPWR _02005_
+ sky130_fd_sc_hd__a21oi_1
X_09536_ _04541_ VGND VGND VPWR VPWR _00071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09467_ _04504_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08418_ u_rf.reg18_q\[12\] _03353_ _03355_ u_rf.reg23_q\[12\] _03609_ VGND VGND VPWR
+ VPWR _03610_ sky130_fd_sc_hd__a221o_1
X_06679_ u_rf.reg0_q\[5\] _01662_ _01568_ u_rf.reg5_q\[5\] VGND VGND VPWR VPWR _01939_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_385 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09398_ u_rf.reg2_q\[15\] _04459_ _04449_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08349_ u_rf.reg18_q\[9\] _03262_ _03263_ u_rf.reg23_q\[9\] _03543_ VGND VGND VPWR
+ VPWR _03544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11360_ _05544_ VGND VGND VPWR VPWR _00892_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10311_ u_decod.rf_ff_res_data_i\[21\] VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__buf_2
XFILLER_0_104_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11291_ u_rf.reg26_q\[28\] u_decod.rf_ff_res_data_i\[28\] _05499_ VGND VGND VPWR
+ VPWR _05508_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10242_ u_decod.rf_ff_res_data_i\[0\] VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__clkbuf_4
X_10173_ _04422_ _04568_ _04825_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12814_ clknet_leaf_7_clk _00851_ net218 VGND VGND VPWR VPWR u_rf.reg26_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12745_ clknet_leaf_22_clk _00782_ net286 VGND VGND VPWR VPWR u_rf.reg24_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12676_ clknet_leaf_105_clk _00713_ net321 VGND VGND VPWR VPWR u_rf.reg22_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11627_ _04776_ u_rf.reg31_q\[26\] _05679_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_219 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11558_ _05649_ VGND VGND VPWR VPWR _00985_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10509_ _04749_ u_rf.reg15_q\[13\] _05089_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11489_ _04774_ u_rf.reg29_q\[25\] _05607_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07720_ u_rf.reg5_q\[26\] _02664_ _02665_ u_rf.reg19_q\[26\] _02937_ VGND VGND VPWR
+ VPWR _02938_ sky130_fd_sc_hd__a221o_1
X_05981_ _01071_ _01253_ VGND VGND VPWR VPWR _01255_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07651_ _02870_ _02871_ _02681_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07582_ u_rf.reg26_q\[23\] _02368_ _01645_ u_rf.reg20_q\[23\] VGND VGND VPWR VPWR
+ _02806_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06602_ u_decod.rs2_data_q\[3\] _01864_ _01497_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09321_ _04408_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_2
X_06533_ u_rf.reg5_q\[2\] _01569_ _01595_ u_rf.reg19_q\[2\] _01798_ VGND VGND VPWR
+ VPWR _01799_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09252_ _04350_ _04356_ _04355_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06464_ u_rf.reg9_q\[1\] _01635_ _01650_ u_rf.reg4_q\[1\] _01731_ VGND VGND VPWR
+ VPWR _01732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09183_ u_decod.pc_q_o\[18\] u_decod.branch_imm_q_o\[18\] VGND VGND VPWR VPWR _04307_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_437 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08203_ u_decod.rf_ff_res_data_i\[2\] _03382_ _03403_ _03404_ VGND VGND VPWR VPWR
+ _03405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06395_ _01512_ _01514_ _01573_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__and3_2
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08134_ _03299_ _03336_ _03337_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08065_ u_rf.reg18_q\[0\] _03262_ _03263_ u_rf.reg23_q\[0\] _03268_ VGND VGND VPWR
+ VPWR _03269_ sky130_fd_sc_hd__a221o_1
X_07016_ u_rf.reg19_q\[12\] _01594_ _01650_ u_rf.reg4_q\[12\] VGND VGND VPWR VPWR
+ _02262_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ _01358_ u_decod.branch_imm_q_o\[21\] u_decod.branch_imm_q_o\[20\] _01363_
+ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__o211a_1
X_07918_ _03126_ _03127_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[30\] sky130_fd_sc_hd__xor2_1
X_08898_ _01297_ u_decod.branch_imm_q_o\[12\] VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__and2_1
X_07849_ u_rf.reg18_q\[29\] _01787_ _02386_ u_rf.reg27_q\[29\] VGND VGND VPWR VPWR
+ _03061_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_3_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10860_ _05279_ VGND VGND VPWR VPWR _00657_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09519_ _04423_ _04531_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_103 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10791_ u_rf.reg19_q\[17\] _04974_ _05235_ VGND VGND VPWR VPWR _05243_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12530_ clknet_leaf_38_clk _00567_ net274 VGND VGND VPWR VPWR u_rf.reg17_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12461_ clknet_leaf_11_clk _00498_ net226 VGND VGND VPWR VPWR u_rf.reg15_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_810 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11412_ _05572_ VGND VGND VPWR VPWR _00916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12392_ clknet_leaf_58_clk _00429_ net291 VGND VGND VPWR VPWR u_rf.reg13_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11343_ _04763_ u_rf.reg27_q\[20\] _05535_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11274_ _05476_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__clkbuf_8
X_10225_ _04926_ VGND VGND VPWR VPWR _00375_ sky130_fd_sc_hd__clkbuf_1
X_13013_ clknet_leaf_74_clk _01050_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[26\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10156_ _04889_ VGND VGND VPWR VPWR _00343_ sky130_fd_sc_hd__clkbuf_1
X_10087_ u_rf.reg9_q\[23\] _04476_ _04849_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10989_ _05348_ VGND VGND VPWR VPWR _00717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12728_ clknet_leaf_68_clk _00765_ net351 VGND VGND VPWR VPWR u_rf.reg23_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12659_ clknet_leaf_68_clk _00696_ net351 VGND VGND VPWR VPWR u_rf.reg21_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_684 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06180_ _01450_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09870_ _04719_ u_rf.reg7_q\[0\] _04722_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03978_ _03985_ _03994_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_55_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ u_rf.reg16_q\[27\] _03450_ _03515_ u_rf.reg5_q\[27\] VGND VGND VPWR VPWR
+ _03929_ sky130_fd_sc_hd__a22o_1
X_05964_ _01234_ _01094_ _01240_ _01242_ VGND VGND VPWR VPWR u_decod.dec0.operation_o\[3\]
+ sky130_fd_sc_hd__a31o_1
X_08683_ u_rf.reg31_q\[24\] _03290_ _03292_ u_rf.reg11_q\[24\] _03862_ VGND VGND VPWR
+ VPWR _03863_ sky130_fd_sc_hd__a221o_1
X_07703_ _02828_ _02921_ _02681_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__mux2_1
X_05895_ net487 _01142_ _01119_ net85 _01188_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__a221o_1
X_07634_ u_rf.reg1_q\[24\] _02604_ _02419_ u_rf.reg28_q\[24\] _02855_ VGND VGND VPWR
+ VPWR _02856_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_812 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07565_ _01481_ _02728_ _02788_ _02789_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09304_ _04397_ u_decod.rs2_data_q\[14\] _04398_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06516_ u_rf.reg29_q\[2\] _01780_ _01639_ u_rf.reg21_q\[2\] _01781_ VGND VGND VPWR
+ VPWR _01782_ sky130_fd_sc_hd__a221o_1
X_07496_ _01425_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09235_ u_decod.pc_q_o\[26\] u_decod.branch_imm_q_o\[26\] VGND VGND VPWR VPWR _04351_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_91_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06447_ _01205_ _01529_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__or2_2
XFILLER_0_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_848 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09166_ _04283_ _04287_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__and2_1
XFILLER_0_44_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06378_ _01512_ _01514_ _01551_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__and3_4
XFILLER_0_142_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09097_ _04231_ _04232_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__and2_1
X_08117_ _03320_ VGND VGND VPWR VPWR _03321_ sky130_fd_sc_hd__buf_6
XFILLER_0_9_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08048_ _03228_ _03252_ _03253_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10010_ _04811_ VGND VGND VPWR VPWR _00275_ sky130_fd_sc_hd__clkbuf_1
X_09999_ u_rf.reg8_q\[14\] _04457_ _04801_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11961_ clknet_leaf_89_clk net470 net360 VGND VGND VPWR VPWR u_decod.pc_q_o\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10912_ _05307_ VGND VGND VPWR VPWR _00681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ clknet_leaf_98_clk u_decod.rs2_data_nxt\[13\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10843_ _05270_ VGND VGND VPWR VPWR _00649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10774_ u_rf.reg19_q\[9\] _04957_ _05224_ VGND VGND VPWR VPWR _05234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12513_ clknet_leaf_16_clk _00550_ net251 VGND VGND VPWR VPWR u_rf.reg17_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_57_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12444_ clknet_leaf_128_clk _00481_ net236 VGND VGND VPWR VPWR u_rf.reg15_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12375_ clknet_leaf_69_clk _00412_ net353 VGND VGND VPWR VPWR u_rf.reg12_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_520 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11326_ _04747_ u_rf.reg27_q\[12\] _05524_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_130_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11257_ _05490_ VGND VGND VPWR VPWR _00843_ sky130_fd_sc_hd__clkbuf_1
X_10208_ _04917_ VGND VGND VPWR VPWR _00367_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_66_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11188_ u_rf.reg25_q\[11\] _04962_ _05452_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__mux2_1
X_10139_ _04880_ VGND VGND VPWR VPWR _00335_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_417 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07350_ net100 net43 _02446_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_75_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06301_ u_rf.reg6_q\[0\] _01557_ _01562_ u_rf.reg7_q\[0\] _01570_ VGND VGND VPWR
+ VPWR _01571_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_415 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09020_ _02621_ _04165_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__nor2_2
X_07281_ u_rf.reg0_q\[17\] _01662_ _01635_ u_rf.reg9_q\[17\] _02516_ VGND VGND VPWR
+ VPWR _02517_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_196 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06232_ _01493_ _01501_ _01502_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06163_ _01433_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06094_ u_decod.rs2_data_q\[20\] _01363_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_84_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09922_ _04757_ u_rf.reg7_q\[17\] _04743_ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__mux2_1
X_09853_ _04712_ VGND VGND VPWR VPWR _00217_ sky130_fd_sc_hd__clkbuf_1
X_09784_ _04675_ VGND VGND VPWR VPWR _00185_ sky130_fd_sc_hd__clkbuf_1
X_08804_ u_rf.reg30_q\[30\] _03341_ _03342_ u_rf.reg10_q\[30\] _03977_ VGND VGND VPWR
+ VPWR _03978_ sky130_fd_sc_hd__a221o_1
X_08735_ _03906_ _03908_ _03910_ _03912_ VGND VGND VPWR VPWR _03913_ sky130_fd_sc_hd__or4_1
X_06996_ net36 _02047_ _02049_ net53 _02051_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05947_ _01071_ u_decod.dec0.funct3\[1\] _01077_ VGND VGND VPWR VPWR _01228_ sky130_fd_sc_hd__a21oi_1
X_08666_ u_rf.reg1_q\[23\] _03446_ _03447_ u_rf.reg14_q\[23\] VGND VGND VPWR VPWR
+ _03847_ sky130_fd_sc_hd__a22o_1
X_05878_ u_exe.pc_data_q\[24\] _01118_ _01100_ net81 VGND VGND VPWR VPWR _01176_ sky130_fd_sc_hd__a22o_1
XANTENNA_108 u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08597_ u_rf.reg9_q\[20\] _03294_ _03296_ u_rf.reg20_q\[20\] _03780_ VGND VGND VPWR
+ VPWR _03781_ sky130_fd_sc_hd__a221o_1
X_07617_ _02334_ _02815_ _02816_ _02839_ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o31a_2
XTAP_TAPCELL_ROW_101_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07548_ u_decod.pc_q_o\[21\] u_decod.pc_q_o\[22\] u_decod.pc_q_o\[23\] _02638_ VGND
+ VGND VPWR VPWR _02773_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_93_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07479_ u_rf.reg16_q\[21\] _01564_ _01630_ u_rf.reg17_q\[21\] VGND VGND VPWR VPWR
+ _02707_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09218_ _04335_ _04336_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__or2b_1
X_10490_ _04730_ u_rf.reg15_q\[4\] _05078_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09149_ _04276_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12160_ clknet_leaf_117_clk _00197_ net323 VGND VGND VPWR VPWR u_rf.reg6_q\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11111_ u_rf.reg24_q\[7\] _04953_ _05405_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12091_ clknet_leaf_11_clk _00128_ net222 VGND VGND VPWR VPWR u_rf.reg4_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11042_ _05376_ VGND VGND VPWR VPWR _00742_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12993_ clknet_leaf_92_clk _01030_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[6\]
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11944_ clknet_leaf_92_clk u_decod.rs1_data_nxt\[32\] net345 VGND VGND VPWR VPWR
+ u_decod.rs1_data_q\[32\] sky130_fd_sc_hd__dfrtp_2
X_11875_ clknet_leaf_98_clk u_decod.dec0.unsign_extension net332 VGND VGND VPWR VPWR
+ u_decod.unsign_ext_q_o sky130_fd_sc_hd__dfrtp_1
X_10826_ u_rf.reg20_q\[1\] _04941_ _05260_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10757_ _05225_ VGND VGND VPWR VPWR _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_768 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_133_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_133_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_124_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10688_ u_rf.reg18_q\[0\] _04935_ _05188_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12427_ clknet_leaf_1_clk _00464_ net221 VGND VGND VPWR VPWR u_rf.reg14_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12358_ clknet_leaf_140_clk _00395_ net204 VGND VGND VPWR VPWR u_rf.reg12_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12289_ clknet_leaf_17_clk _00326_ net251 VGND VGND VPWR VPWR u_rf.reg10_q\[6\] sky130_fd_sc_hd__dfrtp_1
X_11309_ _04730_ u_rf.reg27_q\[4\] _05513_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06850_ _01422_ _02040_ _01441_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05801_ u_decod.pc0_q_i\[6\] net381 VGND VGND VPWR VPWR _01117_ sky130_fd_sc_hd__nand2_1
X_06781_ _01945_ _02036_ net201 VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__a21o_1
X_05732_ _01058_ VGND VGND VPWR VPWR _01059_ sky130_fd_sc_hd__clkbuf_4
X_08520_ _03701_ _03703_ _03705_ _03707_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__or4_1
X_08451_ u_rf.reg0_q\[13\] _03174_ _03291_ u_rf.reg11_q\[13\] VGND VGND VPWR VPWR
+ _03642_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07402_ _02189_ _02585_ _02632_ _01506_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08382_ u_rf.reg15_q\[10\] _03373_ _03374_ u_rf.reg24_q\[10\] _03575_ VGND VGND VPWR
+ VPWR _03576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07333_ u_rf.reg1_q\[18\] _01586_ _01666_ u_rf.reg8_q\[18\] VGND VGND VPWR VPWR _02567_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_63_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_124_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_124_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_34_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07264_ _01475_ _02450_ _02500_ _01478_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__a211o_1
X_09003_ _04149_ _04150_ VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__xor2_1
X_06215_ net98 net99 VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07195_ u_rf.reg23_q\[15\] _01613_ _01622_ u_rf.reg24_q\[15\] VGND VGND VPWR VPWR
+ _02435_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06146_ _01271_ _01416_ _01268_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06077_ u_decod.rs2_data_q\[12\] _01297_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_581 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09905_ _04746_ VGND VGND VPWR VPWR _00235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09836_ _04703_ VGND VGND VPWR VPWR _00209_ sky130_fd_sc_hd__clkbuf_1
X_09767_ _04666_ VGND VGND VPWR VPWR _00177_ sky130_fd_sc_hd__clkbuf_1
X_06979_ _02226_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__inv_2
X_08718_ u_rf.reg18_q\[26\] _03352_ _03354_ u_rf.reg23_q\[26\] VGND VGND VPWR VPWR
+ _03896_ sky130_fd_sc_hd__a22o_1
X_09698_ _04628_ VGND VGND VPWR VPWR _00146_ sky130_fd_sc_hd__clkbuf_1
X_08649_ u_rf.reg1_q\[22\] _03311_ _03333_ u_rf.reg2_q\[22\] _03830_ VGND VGND VPWR
+ VPWR _03831_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11660_ u_decod.dec0.funct7\[3\] _05700_ _02644_ _05704_ VGND VGND VPWR VPWR _01032_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10611_ _05147_ VGND VGND VPWR VPWR _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_115_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_115_clk sky130_fd_sc_hd__clkbuf_16
X_11591_ _04740_ u_rf.reg31_q\[9\] _05657_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10542_ _04782_ u_rf.reg15_q\[29\] _05100_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10473_ _05073_ VGND VGND VPWR VPWR _00476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_497 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ clknet_leaf_31_clk _00249_ net261 VGND VGND VPWR VPWR u_rf.reg7_q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12143_ clknet_leaf_38_clk _00180_ net274 VGND VGND VPWR VPWR u_rf.reg5_q\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12074_ clknet_leaf_29_clk _00111_ net257 VGND VGND VPWR VPWR u_rf.reg3_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_11025_ u_rf.reg22_q\[31\] _05003_ _05332_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ clknet_leaf_43_clk _01013_ net294 VGND VGND VPWR VPWR u_rf.reg31_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11927_ clknet_leaf_87_clk u_decod.rs1_data\[15\] net362 VGND VGND VPWR VPWR u_decod.rs1_data_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11858_ clknet_leaf_35_clk _00085_ net276 VGND VGND VPWR VPWR u_rf.reg0_q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_217 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_19 _01664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11789_ clknet_leaf_83_clk net141 net365 VGND VGND VPWR VPWR u_decod.pc0_q_i\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_10809_ _05252_ VGND VGND VPWR VPWR _00633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_106_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06000_ u_decod.rs2_data_q\[30\] u_decod.rs1_data_q\[30\] VGND VGND VPWR VPWR _01271_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput115 net115 VGND VGND VPWR VPWR adr_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_51_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput104 net104 VGND VGND VPWR VPWR adr_o[12] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_149_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput148 net148 VGND VGND VPWR VPWR icache_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput137 net137 VGND VGND VPWR VPWR icache_adr_o[12] sky130_fd_sc_hd__buf_4
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput126 net126 VGND VGND VPWR VPWR adr_o[3] sky130_fd_sc_hd__buf_2
Xoutput159 net159 VGND VGND VPWR VPWR icache_adr_o[3] sky130_fd_sc_hd__buf_2
X_07951_ u_rf.reg16_q\[31\] _02307_ _02379_ u_rf.reg17_q\[31\] VGND VGND VPWR VPWR
+ _03159_ sky130_fd_sc_hd__a22o_1
X_06902_ _01764_ _02149_ _02150_ _02152_ _01344_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__o32a_1
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07882_ _01477_ _03013_ _03092_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09621_ _04587_ VGND VGND VPWR VPWR _00110_ sky130_fd_sc_hd__clkbuf_1
X_06833_ _02035_ _02036_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__and2b_1
X_09552_ u_rf.reg0_q\[15\] _04459_ _04544_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__mux2_1
X_06764_ u_rf.reg5_q\[7\] _01567_ _01620_ u_rf.reg24_q\[7\] VGND VGND VPWR VPWR _02020_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08503_ u_rf.reg4_q\[16\] _03264_ _03267_ u_rf.reg17_q\[16\] VGND VGND VPWR VPWR
+ _03691_ sky130_fd_sc_hd__a22o_1
X_09483_ u_rf.reg1_q\[15\] _04459_ _04507_ VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06695_ _01442_ _01953_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__nand2_1
X_08434_ u_decod.exe_ff_res_data_i\[12\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[12\]
+ _03625_ VGND VGND VPWR VPWR _03626_ sky130_fd_sc_hd__a221o_2
XFILLER_0_148_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08365_ u_rf.reg27_q\[9\] _03365_ _03320_ u_rf.reg19_q\[9\] VGND VGND VPWR VPWR _03560_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07316_ _02332_ _02533_ _02534_ _02550_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[18\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08296_ u_rf.reg4_q\[6\] _03224_ _03225_ u_rf.reg17_q\[6\] VGND VGND VPWR VPWR _03494_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07247_ u_decod.rf_ff_res_data_i\[16\] _01549_ _01714_ _02465_ _02484_ VGND VGND
+ VPWR VPWR _02485_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_07178_ u_decod.dec0.instr_i\[15\] _01208_ _02256_ VGND VGND VPWR VPWR _02418_ sky130_fd_sc_hd__a21oi_1
X_06129_ u_decod.rs2_data_q\[16\] _01388_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout331 net333 VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_4
Xfanout320 net334 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net354 VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_4
Xfanout342 net343 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__buf_2
Xfanout364 net366 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_4
X_09819_ _04694_ VGND VGND VPWR VPWR _00201_ sky130_fd_sc_hd__clkbuf_1
X_12830_ clknet_leaf_132_clk _00867_ net228 VGND VGND VPWR VPWR u_rf.reg27_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12761_ clknet_leaf_58_clk _00798_ net292 VGND VGND VPWR VPWR u_rf.reg24_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12692_ clknet_leaf_31_clk _00729_ net263 VGND VGND VPWR VPWR u_rf.reg22_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11712_ clknet_leaf_137_clk _00004_ net227 VGND VGND VPWR VPWR u_rf.reg2_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11643_ u_decod.branch_imm_q_o\[1\] _01716_ _05693_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_913 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11574_ _05658_ VGND VGND VPWR VPWR _00992_ sky130_fd_sc_hd__clkbuf_1
Xinput17 icache_instr_i[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
Xinput28 icache_instr_i[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_30_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10525_ _05101_ VGND VGND VPWR VPWR _00500_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_96_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput39 load_data_i[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
X_10456_ _04763_ u_rf.reg14_q\[20\] _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_443 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10387_ _05005_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__buf_6
XFILLER_0_0_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12126_ clknet_leaf_134_clk _00163_ net232 VGND VGND VPWR VPWR u_rf.reg5_q\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_127_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12057_ clknet_leaf_95_clk net440 net327 VGND VGND VPWR VPWR u_decod.rf_ff_rd_adr_q_i\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_144_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11008_ _05358_ VGND VGND VPWR VPWR _00726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_36_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ clknet_leaf_130_clk _00996_ net230 VGND VGND VPWR VPWR u_rf.reg31_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06480_ _01683_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__buf_2
XFILLER_0_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08150_ _03352_ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__buf_8
XFILLER_0_114_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07101_ _01820_ _02343_ _01354_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08081_ _03206_ VGND VGND VPWR VPWR _03285_ sky130_fd_sc_hd__buf_6
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07032_ _01772_ u_decod.exe_ff_res_data_i\[12\] _02277_ VGND VGND VPWR VPWR _02278_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_465 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ _01367_ u_decod.branch_imm_q_o\[23\] _04133_ VGND VGND VPWR VPWR _04134_
+ sky130_fd_sc_hd__a21oi_1
X_07934_ _03133_ _03140_ _03142_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[31\]
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07865_ u_rf.reg30_q\[29\] _01581_ _02364_ u_rf.reg21_q\[29\] _03076_ VGND VGND VPWR
+ VPWR _03077_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09604_ _04578_ VGND VGND VPWR VPWR _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07796_ _03008_ _03010_ _02723_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__mux2_1
X_06816_ u_rf.reg31_q\[8\] _01614_ _01648_ u_rf.reg4_q\[8\] VGND VGND VPWR VPWR _02070_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09535_ u_rf.reg0_q\[7\] _04442_ _04533_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__mux2_1
X_06747_ _01480_ _01999_ _02003_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_149_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06678_ u_rf.reg6_q\[5\] _01555_ _01583_ u_rf.reg11_q\[5\] _01937_ VGND VGND VPWR
+ VPWR _01938_ sky130_fd_sc_hd__a221o_1
X_09466_ u_rf.reg1_q\[7\] _04442_ _04496_ VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08417_ u_rf.reg4_q\[12\] _03356_ _03357_ u_rf.reg17_q\[12\] VGND VGND VPWR VPWR
+ _03609_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_397 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09397_ u_decod.rf_ff_res_data_i\[15\] VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__buf_2
XFILLER_0_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08348_ u_rf.reg4_q\[9\] _03265_ _03267_ u_rf.reg17_q\[9\] VGND VGND VPWR VPWR _03543_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08279_ u_decod.exe_ff_res_data_i\[5\] _03381_ _03477_ VGND VGND VPWR VPWR _03478_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11290_ _05507_ VGND VGND VPWR VPWR _00859_ sky130_fd_sc_hd__clkbuf_1
X_10310_ _04982_ VGND VGND VPWR VPWR _00404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10241_ _04934_ VGND VGND VPWR VPWR _00383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_91_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10172_ _04897_ VGND VGND VPWR VPWR _00351_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12813_ clknet_leaf_7_clk _00850_ net217 VGND VGND VPWR VPWR u_rf.reg26_q\[18\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12744_ clknet_leaf_59_clk _00781_ net290 VGND VGND VPWR VPWR u_rf.reg24_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12675_ clknet_leaf_105_clk _00712_ net320 VGND VGND VPWR VPWR u_rf.reg22_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11626_ _05685_ VGND VGND VPWR VPWR _01017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ _04774_ u_rf.reg30_q\[25\] _05643_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_708 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10508_ _05092_ VGND VGND VPWR VPWR _00492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11488_ _05612_ VGND VGND VPWR VPWR _00952_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10439_ _04747_ u_rf.reg14_q\[12\] _05053_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12109_ clknet_leaf_6_clk _00146_ net215 VGND VGND VPWR VPWR u_rf.reg4_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_05980_ _01254_ VGND VGND VPWR VPWR u_decod.dec0.access_size_o\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07650_ _01472_ _02679_ _01500_ VGND VGND VPWR VPWR _02871_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07581_ u_rf.reg0_q\[23\] _01664_ _02371_ u_rf.reg15_q\[23\] _02804_ VGND VGND VPWR
+ VPWR _02805_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06601_ _01322_ _01494_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__and2_1
X_09320_ _04397_ u_decod.rs2_data_q\[22\] _04398_ VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and3_1
XFILLER_0_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06532_ u_rf.reg16_q\[2\] _01565_ _01631_ u_rf.reg17_q\[2\] VGND VGND VPWR VPWR _01798_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09251_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08202_ _03253_ VGND VGND VPWR VPWR _03404_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06463_ u_rf.reg18_q\[1\] _01591_ _01612_ u_rf.reg23_q\[1\] VGND VGND VPWR VPWR _01731_
+ sky130_fd_sc_hd__a22o_1
X_06394_ _01663_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__buf_6
X_09182_ u_decod.pc_q_o\[18\] u_decod.branch_imm_q_o\[18\] VGND VGND VPWR VPWR _04306_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_90_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08133_ _03253_ VGND VGND VPWR VPWR _03337_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08064_ u_rf.reg4_q\[0\] _03265_ _03267_ u_rf.reg17_q\[0\] VGND VGND VPWR VPWR _03268_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_776 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07015_ u_rf.reg31_q\[12\] _01616_ _01659_ u_rf.reg14_q\[12\] _02260_ VGND VGND VPWR
+ VPWR _02261_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_73_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ _04117_ _04118_ VGND VGND VPWR VPWR _04119_ sky130_fd_sc_hd__nand2_1
X_07917_ _03041_ _03042_ _03081_ _01897_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__o31a_1
X_08897_ _01297_ u_decod.branch_imm_q_o\[12\] VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_95_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_07848_ u_decod.dec0.funct7\[4\] _01224_ _02646_ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07779_ _01528_ _02929_ _02951_ _02953_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_104_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ u_decod.rf_ff_rd_adr_q_i\[0\] _04424_ _01531_ _01536_ VGND VGND VPWR VPWR
+ _04531_ sky130_fd_sc_hd__or4_4
XFILLER_0_78_240 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10790_ _05242_ VGND VGND VPWR VPWR _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09449_ _01534_ _04424_ _01531_ _01536_ VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__or4_4
XFILLER_0_152_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12460_ clknet_leaf_20_clk _00497_ net280 VGND VGND VPWR VPWR u_rf.reg15_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11411_ u_rf.reg28_q\[20\] u_decod.rf_ff_res_data_i\[20\] _05571_ VGND VGND VPWR
+ VPWR _05572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12391_ clknet_leaf_5_clk _00428_ net213 VGND VGND VPWR VPWR u_rf.reg13_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11342_ _05512_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__buf_6
XFILLER_0_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11273_ _05498_ VGND VGND VPWR VPWR _00851_ sky130_fd_sc_hd__clkbuf_1
X_10224_ _04770_ u_rf.reg11_q\[23\] _04922_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__mux2_1
X_13012_ clknet_leaf_74_clk _01049_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[25\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10155_ u_rf.reg10_q\[23\] _04476_ _04885_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10086_ _04852_ VGND VGND VPWR VPWR _00310_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_86_clk clknet_4_11_0_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_113_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10988_ u_rf.reg22_q\[13\] _04966_ _05344_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__mux2_1
X_12727_ clknet_leaf_70_clk _00764_ net352 VGND VGND VPWR VPWR u_rf.reg23_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12658_ clknet_leaf_39_clk _00695_ net279 VGND VGND VPWR VPWR u_rf.reg21_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_833 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11609_ _05676_ VGND VGND VPWR VPWR _01009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
X_12589_ clknet_leaf_5_clk _00626_ net217 VGND VGND VPWR VPWR u_rf.reg19_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03987_ _03989_ _03991_ _03993_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_55_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ u_rf.reg7_q\[27\] _03369_ _03370_ u_rf.reg25_q\[27\] _03927_ VGND VGND VPWR
+ VPWR _03928_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_77_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
X_05963_ _01071_ u_decod.dec0.funct3\[2\] _01241_ VGND VGND VPWR VPWR _01242_ sky130_fd_sc_hd__and3_1
X_05894_ _01186_ _01144_ _01187_ VGND VGND VPWR VPWR _01188_ sky130_fd_sc_hd__and3b_1
XFILLER_0_136_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08682_ u_rf.reg9_q\[24\] _03294_ _03296_ u_rf.reg20_q\[24\] VGND VGND VPWR VPWR
+ _03862_ sky130_fd_sc_hd__a22o_1
X_07702_ _01472_ _02725_ _01500_ VGND VGND VPWR VPWR _02921_ sky130_fd_sc_hd__o21a_1
X_07633_ u_rf.reg16_q\[24\] _02307_ _01610_ u_rf.reg12_q\[24\] VGND VGND VPWR VPWR
+ _02855_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07564_ _02781_ _01430_ u_decod.instr_unit_q\[1\] _01427_ VGND VGND VPWR VPWR _02789_
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_0_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_824 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07495_ _02720_ _02677_ _02721_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__a21oi_1
X_06515_ u_rf.reg14_q\[2\] _01659_ _01671_ u_rf.reg27_q\[2\] VGND VGND VPWR VPWR _01781_
+ sky130_fd_sc_hd__a22o_1
X_09303_ _04399_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09234_ u_decod.pc_q_o\[26\] u_decod.branch_imm_q_o\[26\] VGND VGND VPWR VPWR _04350_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06446_ _01206_ _01530_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__or2_2
X_09165_ _04290_ _04291_ VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__and2b_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08116_ _03247_ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__buf_6
X_06377_ u_rf.reg9_q\[0\] _01636_ _01639_ u_rf.reg21_q\[0\] _01646_ VGND VGND VPWR
+ VPWR _01647_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09096_ u_decod.pc_q_o\[6\] u_decod.branch_imm_q_o\[6\] VGND VGND VPWR VPWR _04232_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_142_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08047_ _03186_ _03196_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__and2_4
XFILLER_0_4_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09998_ _04805_ VGND VGND VPWR VPWR _00269_ sky130_fd_sc_hd__clkbuf_1
X_08949_ _04103_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_68_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_11960_ clknet_leaf_87_clk net465 net362 VGND VGND VPWR VPWR u_decod.pc_q_o\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_10911_ u_rf.reg21_q\[9\] _04957_ _05297_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ clknet_leaf_98_clk u_decod.rs2_data_nxt\[12\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10842_ u_rf.reg20_q\[9\] _04957_ _05260_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10773_ _05233_ VGND VGND VPWR VPWR _00616_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12512_ clknet_leaf_114_clk _00549_ net323 VGND VGND VPWR VPWR u_rf.reg17_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12443_ clknet_leaf_11_clk _00480_ net222 VGND VGND VPWR VPWR u_rf.reg15_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12374_ clknet_leaf_51_clk _00411_ net307 VGND VGND VPWR VPWR u_rf.reg12_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11325_ _05526_ VGND VGND VPWR VPWR _00875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11256_ u_rf.reg26_q\[11\] u_decod.rf_ff_res_data_i\[11\] _05488_ VGND VGND VPWR
+ VPWR _05490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10207_ _04753_ u_rf.reg11_q\[15\] _04911_ VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11187_ _05453_ VGND VGND VPWR VPWR _00810_ sky130_fd_sc_hd__clkbuf_1
X_10138_ u_rf.reg10_q\[15\] _04459_ _04874_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__mux2_1
X_10069_ _04843_ VGND VGND VPWR VPWR _00302_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_59_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_50_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_744 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07280_ u_rf.reg19_q\[17\] _01594_ _01649_ u_rf.reg4_q\[17\] VGND VGND VPWR VPWR
+ _02516_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06300_ u_rf.reg16_q\[0\] _01565_ _01569_ u_rf.reg5_q\[0\] VGND VGND VPWR VPWR _01570_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06231_ _01315_ _01496_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__nand2_2
XFILLER_0_26_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06162_ u_decod.instr_unit_q\[0\] u_decod.instr_operation_q\[3\] _01056_ VGND VGND
+ VPWR VPWR _01433_ sky130_fd_sc_hd__and3_1
XFILLER_0_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06093_ u_decod.rs2_data_q\[20\] _01363_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09921_ u_decod.rf_ff_res_data_i\[17\] VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09852_ u_rf.reg6_q\[25\] _04480_ _04706_ VGND VGND VPWR VPWR _04712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08803_ u_rf.reg26_q\[30\] _03344_ _03345_ u_rf.reg21_q\[30\] VGND VGND VPWR VPWR
+ _03977_ sky130_fd_sc_hd__a22o_1
X_09783_ u_rf.reg5_q\[25\] _04480_ _04669_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__mux2_1
X_08734_ u_rf.reg0_q\[26\] _03420_ _03421_ u_rf.reg12_q\[26\] _03911_ VGND VGND VPWR
+ VPWR _03912_ sky130_fd_sc_hd__a221o_1
X_06995_ _02234_ _02235_ _01442_ _02241_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__a2bb2o_1
X_05946_ _01080_ _01226_ VGND VGND VPWR VPWR _01227_ sky130_fd_sc_hd__and2b_1
X_08665_ u_rf.reg15_q\[23\] _03373_ _03374_ u_rf.reg24_q\[23\] _03845_ VGND VGND VPWR
+ VPWR _03846_ sky130_fd_sc_hd__a221o_1
X_05877_ u_decod.pc0_q_i\[24\] _01171_ VGND VGND VPWR VPWR _01175_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_68_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 u_decod.rs1_data_q\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08596_ u_rf.reg31_q\[20\] _03289_ _03291_ u_rf.reg11_q\[20\] VGND VGND VPWR VPWR
+ _03780_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _01260_ _02825_ _02838_ VGND VGND VPWR VPWR _02839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07547_ _01373_ _02738_ _01370_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07478_ _02701_ _02703_ _02705_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__or3_1
XFILLER_0_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09217_ u_decod.pc_q_o\[23\] u_decod.branch_imm_q_o\[23\] VGND VGND VPWR VPWR _04336_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06429_ _01316_ _01697_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09148_ u_decod.pc_q_o\[13\] u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR _04277_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09079_ _04210_ _04214_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11110_ _05412_ VGND VGND VPWR VPWR _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_112_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12090_ clknet_leaf_60_clk _00127_ net289 VGND VGND VPWR VPWR u_rf.reg3_q\[31\] sky130_fd_sc_hd__dfrtp_1
X_11041_ _04734_ u_rf.reg23_q\[6\] _05369_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__mux2_1
X_12992_ clknet_leaf_92_clk _01029_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11943_ clknet_leaf_87_clk u_decod.rs1_data\[31\] net362 VGND VGND VPWR VPWR u_decod.rs1_data_q\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11874_ clknet_leaf_103_clk u_decod.dec0.jalr net336 VGND VGND VPWR VPWR u_decod.instr_operation_q\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10825_ _05261_ VGND VGND VPWR VPWR _00640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10756_ u_rf.reg19_q\[0\] _04935_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_421 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10687_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__buf_6
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12426_ clknet_leaf_27_clk _00463_ net258 VGND VGND VPWR VPWR u_rf.reg14_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12357_ clknet_leaf_121_clk _00394_ net248 VGND VGND VPWR VPWR u_rf.reg12_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12288_ clknet_leaf_115_clk _00325_ net323 VGND VGND VPWR VPWR u_rf.reg10_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11308_ _05517_ VGND VGND VPWR VPWR _00867_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11239_ u_rf.reg26_q\[3\] net491 _05477_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05800_ u_decod.pc0_q_i\[6\] net381 VGND VGND VPWR VPWR _01116_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06780_ _01944_ _01990_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__nor2_1
X_05731_ _01057_ VGND VGND VPWR VPWR _01058_ sky130_fd_sc_hd__inv_2
X_08450_ u_rf.reg15_q\[13\] _03300_ _03311_ u_rf.reg1_q\[13\] _03640_ VGND VGND VPWR
+ VPWR _03641_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07401_ _01423_ _02631_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__or2_1
X_08381_ u_rf.reg6_q\[10\] _03305_ _03307_ u_rf.reg13_q\[10\] VGND VGND VPWR VPWR
+ _03575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07332_ u_rf.reg20_q\[18\] _01645_ _01671_ u_rf.reg27_q\[18\] _02565_ VGND VGND VPWR
+ VPWR _02566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07263_ _01493_ _02340_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09002_ _04143_ _04145_ _04142_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07194_ u_rf.reg16_q\[15\] _02307_ _01776_ u_rf.reg2_q\[15\] _02433_ VGND VGND VPWR
+ VPWR _02434_ sky130_fd_sc_hd__a221o_1
X_06214_ _01484_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__buf_4
XFILLER_0_54_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06145_ _01272_ _01415_ _01269_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06076_ _01296_ _01295_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09904_ _04745_ u_rf.reg7_q\[11\] _04743_ VGND VGND VPWR VPWR _04746_ sky130_fd_sc_hd__mux2_1
X_09835_ u_rf.reg6_q\[17\] _04463_ _04695_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09766_ u_rf.reg5_q\[17\] _04463_ _04658_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__mux2_1
X_06978_ _02177_ _02178_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__or2_1
X_08717_ net455 _03773_ _03895_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[25\]
+ sky130_fd_sc_hd__a22o_1
X_05929_ net508 u_decod.dec0.rd_v VGND VGND VPWR VPWR _01216_ sky130_fd_sc_hd__and2_1
X_09697_ u_rf.reg4_q\[18\] _04465_ _04619_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__mux2_1
X_08648_ u_rf.reg13_q\[22\] _03306_ _03285_ u_rf.reg21_q\[22\] VGND VGND VPWR VPWR
+ _03830_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08579_ u_rf.reg27_q\[19\] _03318_ _03320_ u_rf.reg19_q\[19\] VGND VGND VPWR VPWR
+ _03764_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10610_ u_rf.reg16_q\[28\] _04997_ _05138_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_544 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11590_ _05666_ VGND VGND VPWR VPWR _01000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10541_ _05109_ VGND VGND VPWR VPWR _00508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10472_ _04780_ u_rf.reg14_q\[28\] _05064_ VGND VGND VPWR VPWR _05073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12211_ clknet_leaf_67_clk _00248_ net349 VGND VGND VPWR VPWR u_rf.reg7_q\[24\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12142_ clknet_leaf_6_clk _00179_ net216 VGND VGND VPWR VPWR u_rf.reg5_q\[19\] sky130_fd_sc_hd__dfrtp_1
X_12073_ clknet_leaf_24_clk _00110_ net265 VGND VGND VPWR VPWR u_rf.reg3_q\[14\] sky130_fd_sc_hd__dfrtp_1
X_11024_ _05366_ VGND VGND VPWR VPWR _00734_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12975_ clknet_leaf_43_clk _01012_ net294 VGND VGND VPWR VPWR u_rf.reg31_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11926_ clknet_leaf_86_clk u_decod.rs1_data\[14\] net362 VGND VGND VPWR VPWR u_decod.rs1_data_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11857_ clknet_leaf_42_clk _00084_ net276 VGND VGND VPWR VPWR u_rf.reg0_q\[20\] sky130_fd_sc_hd__dfrtp_1
X_11788_ clknet_leaf_83_clk net140 net365 VGND VGND VPWR VPWR u_decod.pc0_q_i\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10808_ u_rf.reg19_q\[25\] _04991_ _05246_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10739_ _05215_ VGND VGND VPWR VPWR _00600_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput116 net116 VGND VGND VPWR VPWR adr_o[23] sky130_fd_sc_hd__buf_2
X_12409_ clknet_leaf_61_clk _00446_ net343 VGND VGND VPWR VPWR u_rf.reg13_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput105 net105 VGND VGND VPWR VPWR adr_o[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput138 net138 VGND VGND VPWR VPWR icache_adr_o[13] sky130_fd_sc_hd__buf_4
Xoutput149 net149 VGND VGND VPWR VPWR icache_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput127 net127 VGND VGND VPWR VPWR adr_o[4] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_149_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07950_ u_rf.reg0_q\[31\] _01664_ _02371_ u_rf.reg15_q\[31\] _03157_ VGND VGND VPWR
+ VPWR _03158_ sky130_fd_sc_hd__a221o_1
X_06901_ _01303_ _01763_ _01819_ _02151_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07881_ _02681_ _03091_ VGND VGND VPWR VPWR _03092_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09620_ u_rf.reg3_q\[14\] _04457_ _04582_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__mux2_1
X_06832_ _01895_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__inv_2
X_09551_ _04549_ VGND VGND VPWR VPWR _00078_ sky130_fd_sc_hd__clkbuf_1
X_06763_ u_rf.reg12_q\[7\] _01608_ _01638_ u_rf.reg21_q\[7\] _02018_ VGND VGND VPWR
+ VPWR _02019_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08502_ net462 _03565_ _03690_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09482_ _04512_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06694_ _01911_ _01952_ _01423_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08433_ _03615_ _03624_ _03337_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o21a_2
XFILLER_0_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08364_ u_rf.reg0_q\[9\] _03420_ _03421_ u_rf.reg12_q\[9\] _03558_ VGND VGND VPWR
+ VPWR _03559_ sky130_fd_sc_hd__a221o_1
X_07315_ _01443_ _02537_ _02547_ _02549_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_116_454 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08295_ u_rf.reg8_q\[6\] _03216_ _03272_ u_rf.reg29_q\[6\] _03492_ VGND VGND VPWR
+ VPWR _03493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07246_ _02467_ _02476_ _02483_ _01679_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__o31a_2
XFILLER_0_131_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07177_ _01437_ _02398_ _02415_ _02417_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[15\]
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06128_ u_decod.rs2_data_q\[23\] _01367_ _01397_ _01398_ _01372_ VGND VGND VPWR VPWR
+ _01399_ sky130_fd_sc_hd__o221a_1
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06059_ _01328_ _01329_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout310 net311 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__buf_4
Xfanout332 net333 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_4
Xfanout321 net322 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_4
Xfanout354 net359 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_2
Xfanout365 net366 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__buf_2
Xfanout343 net348 VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_4
X_09818_ u_rf.reg6_q\[9\] _04446_ _04684_ VGND VGND VPWR VPWR _04694_ sky130_fd_sc_hd__mux2_1
X_09749_ u_rf.reg5_q\[9\] _04446_ _04647_ VGND VGND VPWR VPWR _04657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ clknet_leaf_57_clk _00797_ net343 VGND VGND VPWR VPWR u_rf.reg24_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ clknet_leaf_51_clk _00728_ net305 VGND VGND VPWR VPWR u_rf.reg22_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11711_ clknet_leaf_123_clk _00003_ net241 VGND VGND VPWR VPWR u_rf.reg2_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11642_ _05694_ VGND VGND VPWR VPWR _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11573_ _04719_ u_rf.reg31_q\[0\] _05657_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__mux2_1
Xinput18 icache_instr_i[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10524_ _04763_ u_rf.reg15_q\[20\] _05100_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput29 icache_instr_i[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_1
XFILLER_0_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10455_ _05041_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__buf_6
XFILLER_0_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10386_ _05027_ VGND VGND VPWR VPWR _00435_ sky130_fd_sc_hd__clkbuf_1
X_12125_ clknet_leaf_14_clk _00162_ net244 VGND VGND VPWR VPWR u_rf.reg5_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_499 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12056_ clknet_leaf_95_clk net446 net333 VGND VGND VPWR VPWR u_decod.rf_ff_rd_adr_q_i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11007_ u_rf.reg22_q\[22\] _04985_ _05355_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ clknet_leaf_123_clk _00995_ net232 VGND VGND VPWR VPWR u_rf.reg31_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11909_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[30\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[30\] sky130_fd_sc_hd__dfrtp_1
X_12889_ clknet_leaf_64_clk _00926_ net346 VGND VGND VPWR VPWR u_rf.reg28_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_527 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07100_ _01763_ _02244_ _01293_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08080_ _03203_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__buf_8
XFILLER_0_140_232 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07031_ u_decod.rf_ff_res_data_i\[12\] _01550_ _01773_ _02257_ _02276_ VGND VGND
+ VPWR VPWR _02277_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08982_ _01371_ u_decod.branch_imm_q_o\[22\] _04124_ VGND VGND VPWR VPWR _04133_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_11_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07933_ u_decod.pc_q_o\[31\] _03087_ _03141_ VGND VGND VPWR VPWR _03142_ sky130_fd_sc_hd__a21o_1
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07864_ u_rf.reg6_q\[29\] _01557_ _01654_ u_rf.reg22_q\[29\] VGND VGND VPWR VPWR
+ _03076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09603_ u_rf.reg3_q\[6\] _04440_ _04571_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__mux2_1
X_06815_ u_rf.reg29_q\[8\] _01626_ _01637_ u_rf.reg21_q\[8\] _02068_ VGND VGND VPWR
+ VPWR _02069_ sky130_fd_sc_hd__a221o_1
X_07795_ _02921_ _03009_ _02681_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__mux2_1
X_09534_ _04540_ VGND VGND VPWR VPWR _00070_ sky130_fd_sc_hd__clkbuf_1
X_06746_ _01424_ _02002_ _01506_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_628 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09465_ _04503_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
X_06677_ u_rf.reg7_q\[5\] _01560_ _01604_ u_rf.reg3_q\[5\] VGND VGND VPWR VPWR _01937_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_436 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08416_ u_rf.reg8_q\[12\] _03407_ _03408_ u_rf.reg29_q\[12\] _03607_ VGND VGND VPWR
+ VPWR _03608_ sky130_fd_sc_hd__a221o_1
X_09396_ _04458_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_661 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_683 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08347_ net474 _03259_ _03542_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[8\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08278_ u_decod.rf_ff_res_data_i\[5\] _03382_ _03476_ _03404_ VGND VGND VPWR VPWR
+ _03477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07229_ u_rf.reg16_q\[16\] _01565_ _01674_ u_rf.reg2_q\[16\] _02466_ VGND VGND VPWR
+ VPWR _02467_ sky130_fd_sc_hd__a221o_1
X_10240_ _04786_ u_rf.reg11_q\[31\] _04899_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_652 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10171_ u_rf.reg10_q\[31\] _04492_ _04862_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12812_ clknet_leaf_20_clk _00849_ net280 VGND VGND VPWR VPWR u_rf.reg26_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12743_ clknet_leaf_4_clk _00780_ net212 VGND VGND VPWR VPWR u_rf.reg24_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12674_ clknet_leaf_132_clk _00711_ net230 VGND VGND VPWR VPWR u_rf.reg22_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_11625_ _04774_ u_rf.reg31_q\[25\] _05679_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _05648_ VGND VGND VPWR VPWR _00984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_796 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10507_ _04747_ u_rf.reg15_q\[12\] _05089_ VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11487_ _04772_ u_rf.reg29_q\[24\] _05607_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_591 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_764 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10438_ _05055_ VGND VGND VPWR VPWR _00459_ sky130_fd_sc_hd__clkbuf_1
X_10369_ _04745_ u_rf.reg13_q\[11\] _05017_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12108_ clknet_leaf_9_clk _00145_ net226 VGND VGND VPWR VPWR u_rf.reg4_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12039_ clknet_leaf_96_clk u_decod.exe_ff_res_data_i\[19\] net333 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[19\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07580_ u_rf.reg7_q\[23\] _01561_ _01606_ u_rf.reg3_q\[23\] VGND VGND VPWR VPWR _02804_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06600_ _01322_ _01432_ _01859_ _01862_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__a211o_1
X_06531_ u_rf.reg0_q\[2\] _01663_ _01601_ u_rf.reg15_q\[2\] _01796_ VGND VGND VPWR
+ VPWR _01797_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09250_ _04360_ _04363_ _04346_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_157_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08201_ _03384_ _03393_ _03402_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__or3_2
XFILLER_0_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06462_ u_rf.reg19_q\[1\] _01594_ _01658_ u_rf.reg14_q\[1\] _01729_ VGND VGND VPWR
+ VPWR _01730_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09181_ _04093_ _04274_ _04275_ _04305_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[17\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06393_ _01662_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08132_ _03309_ _03317_ _03327_ _03335_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08063_ _03266_ VGND VGND VPWR VPWR _03267_ sky130_fd_sc_hd__buf_6
XFILLER_0_114_722 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07014_ u_rf.reg7_q\[12\] _01560_ _01642_ u_rf.reg26_q\[12\] VGND VGND VPWR VPWR
+ _02260_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08965_ _01371_ u_decod.branch_imm_q_o\[22\] VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__or2_1
X_07916_ _02357_ u_decod.exe_ff_res_data_i\[30\] _03125_ VGND VGND VPWR VPWR _03126_
+ sky130_fd_sc_hd__a21o_1
X_08896_ _04042_ _04059_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__nor2_1
X_07847_ _03059_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[29\] sky130_fd_sc_hd__inv_2
XFILLER_0_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07778_ _02357_ u_decod.exe_ff_res_data_i\[27\] _02993_ VGND VGND VPWR VPWR _02994_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09517_ _04530_ VGND VGND VPWR VPWR _00063_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06729_ _01977_ _01986_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__or2_1
XFILLER_0_149_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_296 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09448_ _04493_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09379_ u_rf.reg2_q\[9\] _04446_ _04428_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__mux2_1
X_11410_ _05548_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12390_ clknet_leaf_139_clk _00427_ net203 VGND VGND VPWR VPWR u_rf.reg13_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_593 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11341_ _05534_ VGND VGND VPWR VPWR _00883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11272_ u_rf.reg26_q\[19\] u_decod.rf_ff_res_data_i\[19\] _05488_ VGND VGND VPWR
+ VPWR _05498_ sky130_fd_sc_hd__mux2_1
X_13011_ clknet_leaf_74_clk _01048_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[24\]
+ sky130_fd_sc_hd__dfxtp_1
X_10223_ _04925_ VGND VGND VPWR VPWR _00374_ sky130_fd_sc_hd__clkbuf_1
X_10154_ _04888_ VGND VGND VPWR VPWR _00342_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10085_ u_rf.reg9_q\[22\] _04474_ _04849_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10987_ _05347_ VGND VGND VPWR VPWR _00716_ sky130_fd_sc_hd__clkbuf_1
X_12726_ clknet_leaf_49_clk _00763_ net309 VGND VGND VPWR VPWR u_rf.reg23_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_139_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_756 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12657_ clknet_leaf_55_clk _00694_ net287 VGND VGND VPWR VPWR u_rf.reg21_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11608_ _04757_ u_rf.reg31_q\[17\] _05668_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ clknet_leaf_26_clk _00625_ net265 VGND VGND VPWR VPWR u_rf.reg19_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_152_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11539_ _05639_ VGND VGND VPWR VPWR _00976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08750_ u_rf.reg1_q\[27\] _03446_ _03447_ u_rf.reg14_q\[27\] VGND VGND VPWR VPWR
+ _03927_ sky130_fd_sc_hd__a22o_1
X_05962_ _01068_ _01201_ VGND VGND VPWR VPWR _01241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05893_ u_decod.pc0_q_i\[26\] u_decod.pc0_q_i\[27\] _01177_ u_decod.pc0_q_i\[28\]
+ VGND VGND VPWR VPWR _01187_ sky130_fd_sc_hd__a31o_1
X_08681_ u_rf.reg30_q\[24\] _03281_ _03283_ u_rf.reg10_q\[24\] _03860_ VGND VGND VPWR
+ VPWR _03861_ sky130_fd_sc_hd__a221o_1
X_07701_ _02875_ _02919_ _01481_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__mux2_1
X_07632_ u_rf.reg0_q\[24\] _01664_ _01787_ u_rf.reg18_q\[24\] _02853_ VGND VGND VPWR
+ VPWR _02854_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07563_ _01480_ _02787_ VGND VGND VPWR VPWR _02788_ sky130_fd_sc_hd__nor2_1
X_09302_ _04397_ u_decod.rs2_data_q\[13\] _04398_ VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07494_ u_decod.pc_q_o\[21\] u_decod.pc_q_o\[22\] _02638_ _02334_ VGND VGND VPWR
+ VPWR _02721_ sky130_fd_sc_hd__a31o_1
X_06514_ _01628_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__buf_6
XFILLER_0_64_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09233_ _04141_ _04206_ _04197_ _04349_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[25\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06445_ _01518_ _01527_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__nor2_4
XFILLER_0_8_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09164_ u_decod.pc_q_o\[15\] u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR _04291_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08115_ _03318_ VGND VGND VPWR VPWR _03319_ sky130_fd_sc_hd__buf_6
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06376_ u_rf.reg26_q\[0\] _01642_ _01645_ u_rf.reg20_q\[0\] VGND VGND VPWR VPWR _01646_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09095_ u_decod.pc_q_o\[6\] u_decod.branch_imm_q_o\[6\] VGND VGND VPWR VPWR _04231_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08046_ _03234_ _03240_ _03245_ _03251_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09997_ u_rf.reg8_q\[13\] _04455_ _04801_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__mux2_1
X_08948_ _04096_ _04099_ _04095_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_4_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08879_ _04043_ _04044_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__nor2_1
X_10910_ _05306_ VGND VGND VPWR VPWR _00680_ sky130_fd_sc_hd__clkbuf_1
X_11890_ clknet_leaf_99_clk u_decod.rs2_data_nxt\[11\] net329 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10841_ _05269_ VGND VGND VPWR VPWR _00648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_553 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10772_ u_rf.reg19_q\[8\] _04955_ _05224_ VGND VGND VPWR VPWR _05233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12511_ clknet_leaf_136_clk _00548_ net205 VGND VGND VPWR VPWR u_rf.reg17_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12442_ clknet_leaf_60_clk _00479_ net340 VGND VGND VPWR VPWR u_rf.reg14_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12373_ clknet_leaf_44_clk _00410_ net296 VGND VGND VPWR VPWR u_rf.reg12_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_686 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11324_ _04745_ u_rf.reg27_q\[11\] _05524_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11255_ _05489_ VGND VGND VPWR VPWR _00842_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10206_ _04916_ VGND VGND VPWR VPWR _00366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11186_ u_rf.reg25_q\[10\] _04959_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__mux2_1
X_10137_ _04879_ VGND VGND VPWR VPWR _00334_ sky130_fd_sc_hd__clkbuf_1
X_10068_ u_rf.reg9_q\[14\] _04457_ _04838_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_358 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_778 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12709_ clknet_leaf_125_clk _00746_ net240 VGND VGND VPWR VPWR u_rf.reg23_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06230_ _01451_ _01499_ _01500_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_86 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06161_ _01431_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__buf_4
X_06092_ u_decod.rs1_data_q\[20\] VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09920_ _04756_ VGND VGND VPWR VPWR _00240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09851_ _04711_ VGND VGND VPWR VPWR _00216_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09782_ _04674_ VGND VGND VPWR VPWR _00184_ sky130_fd_sc_hd__clkbuf_1
X_08802_ net451 _03773_ _03976_ _03794_ VGND VGND VPWR VPWR u_decod.rs1_data\[29\]
+ sky130_fd_sc_hd__a22o_1
X_06994_ _02194_ _02240_ _01423_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ u_rf.reg28_q\[26\] _03556_ _03557_ u_rf.reg2_q\[26\] VGND VGND VPWR VPWR
+ _03911_ sky130_fd_sc_hd__a22o_1
X_05945_ u_decod.dec0.instr_i\[4\] _01225_ VGND VGND VPWR VPWR _01226_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08664_ u_rf.reg6_q\[23\] _03304_ _03307_ u_rf.reg13_q\[23\] VGND VGND VPWR VPWR
+ _03845_ sky130_fd_sc_hd__a22o_1
X_05876_ u_decod.pc0_q_i\[24\] _01171_ VGND VGND VPWR VPWR _01174_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_818 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08595_ u_rf.reg30_q\[20\] _03281_ _03283_ u_rf.reg10_q\[20\] _03778_ VGND VGND VPWR
+ VPWR _03779_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ _01443_ _02826_ _02831_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07546_ _01398_ _02770_ _02738_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__or3b_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_715 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09216_ u_decod.pc_q_o\[23\] u_decod.branch_imm_q_o\[23\] VGND VGND VPWR VPWR _04335_
+ sky130_fd_sc_hd__nor2_1
X_07477_ u_rf.reg13_q\[21\] _01598_ _01592_ u_rf.reg18_q\[21\] _02704_ VGND VGND VPWR
+ VPWR _02705_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06428_ u_decod.instr_operation_q\[3\] _01259_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__nand2_2
XFILLER_0_9_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09147_ u_decod.pc_q_o\[13\] u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR _04276_
+ sky130_fd_sc_hd__nor2_1
X_06359_ _01538_ _01515_ _01566_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__and3_4
XFILLER_0_44_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_121_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09078_ _04215_ _04216_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08029_ _03171_ _03199_ _03205_ VGND VGND VPWR VPWR _03235_ sky130_fd_sc_hd__and3_4
XFILLER_0_31_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_141_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11040_ _05375_ VGND VGND VPWR VPWR _00741_ sky130_fd_sc_hd__clkbuf_1
X_12991_ clknet_leaf_93_clk _01028_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[4\]
+ sky130_fd_sc_hd__dfxtp_2
X_11942_ clknet_leaf_65_clk u_decod.rs1_data\[30\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_28_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ clknet_leaf_104_clk u_decod.dec0.operation_o\[4\] net335 VGND VGND VPWR VPWR
+ u_decod.instr_operation_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10824_ u_rf.reg20_q\[0\] _04935_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10755_ _05223_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__buf_6
XFILLER_0_27_428 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_433 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10686_ _04426_ _05114_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__nor2_4
X_12425_ clknet_leaf_19_clk _00462_ net282 VGND VGND VPWR VPWR u_rf.reg14_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12356_ clknet_leaf_112_clk _00393_ net317 VGND VGND VPWR VPWR u_rf.reg12_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11307_ _04728_ u_rf.reg27_q\[3\] _05513_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12287_ clknet_leaf_131_clk _00324_ net227 VGND VGND VPWR VPWR u_rf.reg10_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11238_ _05480_ VGND VGND VPWR VPWR _00834_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11169_ u_rf.reg25_q\[2\] _04943_ _05441_ VGND VGND VPWR VPWR _05444_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_05730_ u_decod.instr_unit_q\[3\] _01056_ VGND VGND VPWR VPWR _01057_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07400_ _02541_ _02630_ _01475_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08380_ _03567_ _03569_ _03571_ _03573_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__or4_1
XFILLER_0_86_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07331_ u_rf.reg23_q\[18\] _01613_ _01622_ u_rf.reg24_q\[18\] VGND VGND VPWR VPWR
+ _02565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07262_ _02197_ _02294_ _02400_ _02498_ _01474_ _01905_ VGND VGND VPWR VPWR _02499_
+ sky130_fd_sc_hd__mux4_2
XTAP_TAPCELL_ROW_14_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09001_ _04147_ _04148_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07193_ u_rf.reg1_q\[15\] _01587_ _01667_ u_rf.reg8_q\[15\] VGND VGND VPWR VPWR _02433_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06213_ _01483_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_680 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06144_ _01262_ _01264_ _01414_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_308 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06075_ _01305_ _01308_ _01341_ _01342_ _01345_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__o311a_1
XFILLER_0_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09903_ u_decod.rf_ff_res_data_i\[11\] VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _04702_ VGND VGND VPWR VPWR _00208_ sky130_fd_sc_hd__clkbuf_1
X_06977_ _01772_ u_decod.exe_ff_res_data_i\[11\] _02224_ VGND VGND VPWR VPWR _02225_
+ sky130_fd_sc_hd__a21o_1
X_09765_ _04665_ VGND VGND VPWR VPWR _00176_ sky130_fd_sc_hd__clkbuf_1
X_08716_ u_decod.exe_ff_res_data_i\[25\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[25\]
+ _03894_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__a221o_1
Xrebuffer30 _01129_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_1
X_09696_ _04627_ VGND VGND VPWR VPWR _00145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_05928_ _01215_ VGND VGND VPWR VPWR u_decod.dec0.rd_o\[1\] sky130_fd_sc_hd__clkbuf_1
X_05859_ net489 _01142_ _01132_ net75 _01161_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__a221o_1
X_08647_ u_rf.reg27_q\[22\] _03318_ _03277_ u_rf.reg3_q\[22\] _03828_ VGND VGND VPWR
+ VPWR _03829_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_83_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08578_ _03756_ _03758_ _03760_ _03762_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__or4_1
XFILLER_0_77_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07529_ u_rf.reg9_q\[22\] _02360_ _02364_ u_rf.reg21_q\[22\] _02754_ VGND VGND VPWR
+ VPWR _02755_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10540_ _04780_ u_rf.reg15_q\[28\] _05100_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_556 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10471_ _05072_ VGND VGND VPWR VPWR _00475_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_98_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_921 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12210_ clknet_leaf_39_clk _00247_ net277 VGND VGND VPWR VPWR u_rf.reg7_q\[23\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_114_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12141_ clknet_leaf_6_clk _00178_ net215 VGND VGND VPWR VPWR u_rf.reg5_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_374 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12072_ clknet_leaf_17_clk _00109_ net288 VGND VGND VPWR VPWR u_rf.reg3_q\[13\] sky130_fd_sc_hd__dfrtp_1
X_11023_ u_rf.reg22_q\[30\] _05001_ _05332_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12974_ clknet_leaf_27_clk _01011_ net258 VGND VGND VPWR VPWR u_rf.reg31_q\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11925_ clknet_leaf_87_clk u_decod.rs1_data\[13\] net360 VGND VGND VPWR VPWR u_decod.rs1_data_q\[13\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_142_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11856_ clknet_leaf_28_clk _00083_ net256 VGND VGND VPWR VPWR u_rf.reg0_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10807_ _05251_ VGND VGND VPWR VPWR _00632_ sky130_fd_sc_hd__clkbuf_1
X_11787_ clknet_leaf_83_clk net139 net365 VGND VGND VPWR VPWR u_decod.pc0_q_i\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10738_ u_rf.reg18_q\[24\] _04989_ _05210_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10669_ _05178_ VGND VGND VPWR VPWR _00567_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ clknet_leaf_52_clk _00445_ net304 VGND VGND VPWR VPWR u_rf.reg13_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput106 net106 VGND VGND VPWR VPWR adr_o[14] sky130_fd_sc_hd__buf_4
XFILLER_0_23_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput117 net117 VGND VGND VPWR VPWR adr_o[24] sky130_fd_sc_hd__buf_2
X_12339_ clknet_leaf_51_clk _00376_ net304 VGND VGND VPWR VPWR u_rf.reg11_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput139 net139 VGND VGND VPWR VPWR icache_adr_o[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_105_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput128 net128 VGND VGND VPWR VPWR adr_o[5] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_149_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06900_ _01303_ _01434_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__nand2_1
X_07880_ _02917_ _03090_ _02685_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__mux2_1
X_06831_ _01093_ _01090_ _01896_ _01079_ _01237_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_37_74 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09550_ u_rf.reg0_q\[14\] _04457_ _04544_ VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__mux2_1
X_06762_ u_rf.reg25_q\[7\] _01574_ _01614_ u_rf.reg31_q\[7\] VGND VGND VPWR VPWR _02018_
+ sky130_fd_sc_hd__a22o_1
X_08501_ u_decod.exe_ff_res_data_i\[15\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[15\]
+ _03689_ VGND VGND VPWR VPWR _03690_ sky130_fd_sc_hd__a221o_1
X_09481_ u_rf.reg1_q\[14\] _04457_ _04507_ VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08432_ _03617_ _03619_ _03621_ _03623_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__or4_1
X_06693_ _01869_ _01951_ _01688_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08363_ u_rf.reg28_q\[9\] _03556_ _03557_ u_rf.reg2_q\[9\] VGND VGND VPWR VPWR _03558_
+ sky130_fd_sc_hd__a22o_1
X_07314_ u_decod.pc_q_o\[18\] _02506_ _02548_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__o21a_1
X_08294_ u_rf.reg22_q\[6\] _03218_ _03219_ u_rf.reg3_q\[6\] VGND VGND VPWR VPWR _03492_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07245_ _02478_ _02480_ _02482_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__or3_1
XFILLER_0_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07176_ u_decod.pc_q_o\[15\] _02335_ _02416_ VGND VGND VPWR VPWR _02417_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06127_ u_decod.rs2_data_q\[22\] _01371_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_93_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_70 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06058_ u_decod.rs2_data_q\[6\] u_decod.rs1_data_q\[6\] VGND VGND VPWR VPWR _01329_
+ sky130_fd_sc_hd__and2_1
Xfanout300 net301 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_4
Xfanout311 net374 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout322 net334 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_4
Xfanout355 net358 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_4
Xfanout366 net367 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_4
Xfanout344 net348 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_4
Xfanout333 net334 VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_4
X_09817_ _04693_ VGND VGND VPWR VPWR _00200_ sky130_fd_sc_hd__clkbuf_1
X_09748_ _04656_ VGND VGND VPWR VPWR _00168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_401 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11710_ clknet_leaf_13_clk _00002_ net245 VGND VGND VPWR VPWR u_rf.reg2_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_09679_ _04618_ VGND VGND VPWR VPWR _00137_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_38_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ clknet_leaf_39_clk _00727_ net278 VGND VGND VPWR VPWR u_rf.reg22_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11641_ u_decod.branch_imm_q_o\[0\] _05692_ _05693_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11572_ _05656_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__buf_6
XFILLER_0_65_876 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10523_ _05077_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__buf_6
XFILLER_0_80_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 icache_instr_i[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10454_ _05063_ VGND VGND VPWR VPWR _00467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10385_ _04761_ u_rf.reg13_q\[19\] _05017_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12124_ clknet_leaf_128_clk _00161_ net236 VGND VGND VPWR VPWR u_rf.reg5_q\[1\] sky130_fd_sc_hd__dfrtp_1
X_12055_ clknet_leaf_95_clk net449 net325 VGND VGND VPWR VPWR u_decod.rf_ff_rd_adr_q_i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11006_ _05357_ VGND VGND VPWR VPWR _00725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12957_ clknet_leaf_15_clk _00994_ net246 VGND VGND VPWR VPWR u_rf.reg31_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12888_ clknet_leaf_66_clk _00925_ net355 VGND VGND VPWR VPWR u_rf.reg28_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_11908_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[29\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11839_ clknet_leaf_13_clk _00066_ net241 VGND VGND VPWR VPWR u_rf.reg0_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_377 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_155_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07030_ _02266_ _02275_ _01679_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__o21a_2
XFILLER_0_140_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08981_ _04131_ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07932_ u_decod.pc_q_o\[31\] _03087_ _01485_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__o21ai_1
X_07863_ u_rf.reg11_q\[29\] _02375_ _02665_ u_rf.reg19_q\[29\] _03074_ VGND VGND VPWR
+ VPWR _03075_ sky130_fd_sc_hd__a221o_1
X_09602_ _04577_ VGND VGND VPWR VPWR _00101_ sky130_fd_sc_hd__clkbuf_1
X_06814_ u_rf.reg14_q\[8\] _01657_ _01669_ u_rf.reg27_q\[8\] VGND VGND VPWR VPWR _02068_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07794_ _01500_ _02827_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__and2_1
X_09533_ u_rf.reg0_q\[6\] _04440_ _04533_ VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06745_ _01705_ _01824_ _01904_ _02001_ _01474_ _01457_ VGND VGND VPWR VPWR _02002_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09464_ u_rf.reg1_q\[6\] _04440_ _04496_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__mux2_1
X_06676_ u_rf.reg17_q\[5\] _01630_ _01644_ u_rf.reg20_q\[5\] _01935_ VGND VGND VPWR
+ VPWR _01936_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09395_ u_rf.reg2_q\[14\] _04457_ _04449_ VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__mux2_1
X_08415_ u_rf.reg22_q\[12\] _03409_ _03410_ u_rf.reg3_q\[12\] VGND VGND VPWR VPWR
+ _03607_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_331 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08346_ u_decod.exe_ff_res_data_i\[8\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[8\]
+ _03541_ VGND VGND VPWR VPWR _03542_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08277_ _03466_ _03475_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07228_ u_rf.reg1_q\[16\] _01587_ _01667_ u_rf.reg8_q\[16\] VGND VGND VPWR VPWR _02466_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07159_ _01467_ _02000_ _02399_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10170_ _04896_ VGND VGND VPWR VPWR _00350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_664 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_710 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12811_ clknet_leaf_11_clk _00848_ net222 VGND VGND VPWR VPWR u_rf.reg26_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12742_ clknet_leaf_139_clk _00779_ net203 VGND VGND VPWR VPWR u_rf.reg24_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12673_ clknet_leaf_16_clk _00710_ net251 VGND VGND VPWR VPWR u_rf.reg22_q\[6\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11624_ _05684_ VGND VGND VPWR VPWR _01016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_651 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11555_ _04772_ u_rf.reg30_q\[24\] _05643_ VGND VGND VPWR VPWR _05648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11486_ _05611_ VGND VGND VPWR VPWR _00951_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10506_ _05091_ VGND VGND VPWR VPWR _00491_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10437_ _04745_ u_rf.reg14_q\[11\] _05053_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10368_ _05018_ VGND VGND VPWR VPWR _00426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10299_ net524 _04974_ _04960_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__mux2_1
X_12107_ clknet_leaf_135_clk _00144_ net208 VGND VGND VPWR VPWR u_rf.reg4_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12038_ clknet_leaf_95_clk u_decod.exe_ff_res_data_i\[18\] net331 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06530_ u_rf.reg7_q\[2\] _01561_ _01606_ u_rf.reg3_q\[2\] VGND VGND VPWR VPWR _01796_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_798 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06461_ u_rf.reg7_q\[1\] _01560_ _01605_ u_rf.reg3_q\[1\] VGND VGND VPWR VPWR _01729_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08200_ _03395_ _03397_ _03399_ _03401_ VGND VGND VPWR VPWR _03402_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09180_ _04302_ _04304_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_407 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06392_ _01516_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08131_ u_rf.reg0_q\[0\] _03176_ _03329_ u_rf.reg12_q\[0\] _03334_ VGND VGND VPWR
+ VPWR _03335_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_734 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08062_ _03225_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__buf_6
XFILLER_0_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07013_ u_rf.reg15_q\[12\] _01601_ _01609_ u_rf.reg12_q\[12\] _02258_ VGND VGND VPWR
+ VPWR _02259_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08964_ _01371_ u_decod.branch_imm_q_o\[22\] VGND VGND VPWR VPWR _04117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07915_ u_decod.rf_ff_res_data_i\[30\] _02358_ _02743_ _03105_ _03124_ VGND VGND
+ VPWR VPWR _03125_ sky130_fd_sc_hd__a221o_1
X_08895_ _04057_ _04058_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__xnor2_1
X_07846_ _02332_ _03045_ _03058_ VGND VGND VPWR VPWR _03059_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07777_ u_decod.rf_ff_res_data_i\[27\] _02358_ _02743_ _02973_ _02992_ VGND VGND
+ VPWR VPWR _02993_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_104_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09516_ u_rf.reg1_q\[31\] _04492_ _04495_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06728_ _01979_ _01981_ _01983_ _01985_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__or4_1
XFILLER_0_149_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09447_ u_rf.reg2_q\[31\] _04492_ _04427_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06659_ _01309_ _01819_ _01697_ _01311_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09378_ u_decod.rf_ff_res_data_i\[9\] VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08329_ u_rf.reg22_q\[8\] _03275_ _03277_ u_rf.reg3_q\[8\] VGND VGND VPWR VPWR _03525_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11340_ _04761_ u_rf.reg27_q\[19\] _05524_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_13010_ clknet_leaf_74_clk _01047_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[23\]
+ sky130_fd_sc_hd__dfxtp_1
X_11271_ _05497_ VGND VGND VPWR VPWR _00850_ sky130_fd_sc_hd__clkbuf_1
X_10222_ _04768_ u_rf.reg11_q\[22\] _04922_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_18_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10153_ u_rf.reg10_q\[22\] _04474_ _04885_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10084_ _04851_ VGND VGND VPWR VPWR _00309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10986_ u_rf.reg22_q\[12\] _04964_ _05344_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__mux2_1
X_12725_ clknet_leaf_44_clk _00762_ net295 VGND VGND VPWR VPWR u_rf.reg23_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ clknet_leaf_36_clk _00693_ net271 VGND VGND VPWR VPWR u_rf.reg21_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11607_ _05675_ VGND VGND VPWR VPWR _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12587_ clknet_leaf_0_clk _00624_ net208 VGND VGND VPWR VPWR u_rf.reg19_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_518 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11538_ _04755_ u_rf.reg30_q\[16\] _05632_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11469_ _05602_ VGND VGND VPWR VPWR _00943_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_48 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07700_ _02834_ _02918_ _01477_ VGND VGND VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
X_05961_ _01075_ _01084_ _01239_ VGND VGND VPWR VPWR _01240_ sky130_fd_sc_hd__a21o_1
X_05892_ u_decod.pc0_q_i\[27\] u_decod.pc0_q_i\[28\] _01180_ VGND VGND VPWR VPWR _01186_
+ sky130_fd_sc_hd__and3_1
X_08680_ u_rf.reg26_q\[24\] _03343_ _03285_ u_rf.reg21_q\[24\] VGND VGND VPWR VPWR
+ _03860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07631_ u_rf.reg31_q\[24\] _01616_ _02380_ u_rf.reg10_q\[24\] VGND VGND VPWR VPWR
+ _02853_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07562_ _02680_ _02786_ _02681_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_724 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09301_ _01427_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__clkbuf_2
X_06513_ u_rf.reg12_q\[2\] _01610_ _01776_ u_rf.reg2_q\[2\] _01778_ VGND VGND VPWR
+ VPWR _01779_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07493_ u_decod.pc_q_o\[22\] VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09232_ _04347_ _04348_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06444_ _01712_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[1\] sky130_fd_sc_hd__buf_1
XFILLER_0_134_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06375_ _01644_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__buf_8
X_09163_ u_decod.pc_q_o\[15\] u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR _04290_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08114_ _03246_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__buf_6
XFILLER_0_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09094_ _04022_ _04207_ _04208_ _04230_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[5\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_114_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08045_ u_rf.reg27_q\[31\] _03246_ _03247_ u_rf.reg19_q\[31\] _03250_ VGND VGND VPWR
+ VPWR _03251_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ _04804_ VGND VGND VPWR VPWR _00268_ sky130_fd_sc_hd__clkbuf_1
X_08947_ _04102_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08878_ u_decod.rs1_data_q\[9\] u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _04044_
+ sky130_fd_sc_hd__and2_1
X_07829_ _01897_ _03042_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10840_ u_rf.reg20_q\[8\] _04955_ _05260_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10771_ _05232_ VGND VGND VPWR VPWR _00615_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12510_ clknet_leaf_1_clk _00547_ net209 VGND VGND VPWR VPWR u_rf.reg17_q\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12441_ clknet_leaf_58_clk _00478_ net292 VGND VGND VPWR VPWR u_rf.reg14_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12372_ clknet_leaf_24_clk _00409_ net269 VGND VGND VPWR VPWR u_rf.reg12_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_698 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
X_11323_ _05525_ VGND VGND VPWR VPWR _00874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11254_ u_rf.reg26_q\[10\] u_decod.rf_ff_res_data_i\[10\] _05488_ VGND VGND VPWR
+ VPWR _05489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_871 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10205_ _04751_ u_rf.reg11_q\[14\] _04911_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__mux2_1
X_11185_ _05440_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__buf_6
XFILLER_0_100_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10136_ u_rf.reg10_q\[14\] _04457_ _04874_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__mux2_1
X_10067_ _04842_ VGND VGND VPWR VPWR _00301_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10969_ u_rf.reg22_q\[4\] _04947_ _05333_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_136_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_136_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12708_ clknet_leaf_107_clk _00745_ net315 VGND VGND VPWR VPWR u_rf.reg23_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12639_ clknet_leaf_132_clk _00676_ net228 VGND VGND VPWR VPWR u_rf.reg21_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06160_ u_decod.instr_unit_q\[0\] _01430_ _01427_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__and3_2
X_06091_ _01361_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_370 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09850_ u_rf.reg6_q\[24\] _04478_ _04706_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__mux2_1
X_09781_ u_rf.reg5_q\[24\] _04478_ _04669_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__mux2_1
X_08801_ u_decod.exe_ff_res_data_i\[29\] _03381_ _03975_ VGND VGND VPWR VPWR _03976_
+ sky130_fd_sc_hd__a21o_1
X_06993_ _02138_ _02239_ _01493_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__mux2_1
X_08732_ u_rf.reg27_q\[26\] _03365_ _03366_ u_rf.reg19_q\[26\] _03909_ VGND VGND VPWR
+ VPWR _03910_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_53_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05944_ u_decod.dec0.instr_i\[5\] _01199_ VGND VGND VPWR VPWR _01225_ sky130_fd_sc_hd__nand2_2
X_08663_ _03837_ _03839_ _03841_ _03843_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__or4_1
X_05875_ net495 _01142_ _01132_ net80 _01173_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__a221o_1
XFILLER_0_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08594_ u_rf.reg26_q\[20\] _03343_ _03286_ u_rf.reg21_q\[20\] VGND VGND VPWR VPWR
+ _03778_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_101_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07614_ net133 _02832_ _02836_ _01746_ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_68_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07545_ _01368_ _01369_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_127_clk clknet_4_2_0_clk VGND VGND VPWR VPWR clknet_leaf_127_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07476_ u_rf.reg23_q\[21\] _01613_ _01791_ u_rf.reg10_q\[21\] VGND VGND VPWR VPWR
+ _02704_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09215_ _04197_ _04331_ _04333_ _04334_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[22\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06427_ u_decod.rs1_data_q\[1\] _01493_ _01431_ VGND VGND VPWR VPWR _01696_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_62_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09146_ _04196_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06358_ _01627_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09077_ u_decod.pc_q_o\[3\] u_decod.branch_imm_q_o\[3\] VGND VGND VPWR VPWR _04216_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06289_ _01512_ _01551_ _01558_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__and3_2
XFILLER_0_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08028_ u_rf.reg7_q\[31\] _03229_ _03230_ u_rf.reg25_q\[31\] _03233_ VGND VGND VPWR
+ VPWR _03234_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09979_ _04795_ VGND VGND VPWR VPWR _00260_ sky130_fd_sc_hd__clkbuf_1
X_12990_ clknet_leaf_93_clk _01027_ VGND VGND VPWR VPWR u_decod.branch_imm_q_o\[3\]
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_28_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ clknet_leaf_75_clk u_decod.rs1_data\[29\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[29\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_679 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11872_ clknet_leaf_103_clk u_decod.dec0.operation_o\[3\] net335 VGND VGND VPWR VPWR
+ u_decod.instr_operation_q\[3\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10823_ _05259_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_118_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_118_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_464 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10754_ _04569_ _05114_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__nor2_4
XFILLER_0_54_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_790 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10685_ _05186_ VGND VGND VPWR VPWR _00575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_568 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_445 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12424_ clknet_leaf_60_clk _00461_ net289 VGND VGND VPWR VPWR u_rf.reg14_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_361 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12355_ clknet_leaf_109_clk _00392_ net314 VGND VGND VPWR VPWR u_rf.reg12_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11306_ _05516_ VGND VGND VPWR VPWR _00866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12286_ clknet_leaf_123_clk _00323_ net231 VGND VGND VPWR VPWR u_rf.reg10_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11237_ u_rf.reg26_q\[2\] net504 _05477_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _05443_ VGND VGND VPWR VPWR _00801_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ u_rf.reg10_q\[6\] _04440_ _04863_ VGND VGND VPWR VPWR _04870_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11099_ u_rf.reg24_q\[1\] _04941_ _05405_ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_307 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_852 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_109_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_109_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07330_ u_rf.reg11_q\[18\] _01584_ _01598_ u_rf.reg13_q\[18\] _02563_ VGND VGND VPWR
+ VPWR _02564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_261 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09000_ u_decod.rs1_data_q\[27\] u_decod.branch_imm_q_o\[27\] VGND VGND VPWR VPWR
+ _04148_ sky130_fd_sc_hd__nand2_1
X_07261_ _01380_ u_decod.rs1_data_q\[9\] net376 _01747_ _01460_ _01461_ VGND VGND
+ VPWR VPWR _02498_ sky130_fd_sc_hd__mux4_2
XFILLER_0_45_259 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07192_ u_rf.reg17_q\[15\] _02379_ _02380_ u_rf.reg10_q\[15\] _02431_ VGND VGND VPWR
+ VPWR _02432_ sky130_fd_sc_hd__a221o_1
X_06212_ u_decod.instr_unit_q\[2\] _01056_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__and2_1
X_06143_ u_decod.rs2_data_q\[29\] u_decod.rs1_data_q\[29\] VGND VGND VPWR VPWR _01414_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_81_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_292 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06074_ _01343_ _01344_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09902_ _04744_ VGND VGND VPWR VPWR _00234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09833_ u_rf.reg6_q\[16\] _04461_ _04695_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__mux2_1
X_06976_ u_decod.rf_ff_res_data_i\[11\] _01550_ _01773_ _02204_ _02223_ VGND VGND
+ VPWR VPWR _02224_ sky130_fd_sc_hd__a221o_1
X_09764_ u_rf.reg5_q\[16\] _04461_ _04658_ VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__mux2_1
X_08715_ _03884_ _03893_ _03378_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__o21a_1
Xrebuffer20 net395 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
X_09695_ u_rf.reg4_q\[17\] _04463_ _04619_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__mux2_1
X_05927_ net511 u_decod.dec0.rd_v VGND VGND VPWR VPWR _01215_ sky130_fd_sc_hd__and2_1
X_05858_ _01159_ _01144_ _01160_ VGND VGND VPWR VPWR _01161_ sky130_fd_sc_hd__and3b_1
X_08646_ u_rf.reg31_q\[22\] _03289_ _03324_ u_rf.reg5_q\[22\] VGND VGND VPWR VPWR
+ _03828_ sky130_fd_sc_hd__a22o_1
Xrebuffer31 _01139_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05789_ net390 u_decod.pc0_q_i\[3\] _01098_ VGND VGND VPWR VPWR _01108_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_92_800 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08577_ u_rf.reg30_q\[19\] _03280_ _03282_ u_rf.reg10_q\[19\] _03761_ VGND VGND VPWR
+ VPWR _03762_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07528_ u_rf.reg12_q\[22\] _01609_ _01674_ u_rf.reg2_q\[22\] VGND VGND VPWR VPWR
+ _02754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07459_ u_decod.rs2_data_q\[21\] _01358_ u_decod.instr_operation_q\[1\] VGND VGND
+ VPWR VPWR _02688_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10470_ _04778_ u_rf.reg14_q\[27\] _05064_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ _04258_ _04260_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12140_ clknet_leaf_26_clk _00177_ net266 VGND VGND VPWR VPWR u_rf.reg5_q\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12071_ clknet_leaf_3_clk _00108_ net211 VGND VGND VPWR VPWR u_rf.reg3_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_11022_ _05365_ VGND VGND VPWR VPWR _00733_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12973_ clknet_leaf_10_clk _01010_ net224 VGND VGND VPWR VPWR u_rf.reg31_q\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11924_ clknet_leaf_86_clk u_decod.rs1_data\[12\] net362 VGND VGND VPWR VPWR u_decod.rs1_data_q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11855_ clknet_leaf_6_clk _00082_ net215 VGND VGND VPWR VPWR u_rf.reg0_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_10806_ u_rf.reg19_q\[24\] _04989_ _05246_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_902 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11786_ clknet_leaf_84_clk net138 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_682 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10737_ _05214_ VGND VGND VPWR VPWR _00599_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_294 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12407_ clknet_leaf_49_clk _00444_ net352 VGND VGND VPWR VPWR u_rf.reg13_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10668_ u_rf.reg17_q\[23\] _04987_ _05174_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10599_ _05141_ VGND VGND VPWR VPWR _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput107 net107 VGND VGND VPWR VPWR adr_o[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_476 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput118 net118 VGND VGND VPWR VPWR adr_o[25] sky130_fd_sc_hd__buf_4
X_12338_ clknet_leaf_40_clk _00375_ net298 VGND VGND VPWR VPWR u_rf.reg11_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput129 net129 VGND VGND VPWR VPWR adr_o[6] sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_149_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12269_ clknet_leaf_4_clk _00306_ net215 VGND VGND VPWR VPWR u_rf.reg9_q\[18\] sky130_fd_sc_hd__dfrtp_1
X_06830_ _01713_ u_decod.exe_ff_res_data_i\[8\] _02083_ VGND VGND VPWR VPWR _02084_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06761_ u_rf.reg14_q\[7\] _01657_ _01649_ u_rf.reg4_q\[7\] _02016_ VGND VGND VPWR
+ VPWR _02017_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08500_ _03679_ _03688_ _03337_ VGND VGND VPWR VPWR _03689_ sky130_fd_sc_hd__o21a_2
X_09480_ _04511_ VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__clkbuf_1
X_06692_ _01949_ _01752_ _01950_ _01754_ _01457_ _01460_ VGND VGND VPWR VPWR _01951_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_144_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08431_ u_rf.reg0_q\[12\] _03176_ _03329_ u_rf.reg12_q\[12\] _03622_ VGND VGND VPWR
+ VPWR _03623_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08362_ _03332_ VGND VGND VPWR VPWR _03557_ sky130_fd_sc_hd__buf_6
XFILLER_0_156_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07313_ u_decod.pc_q_o\[18\] _02506_ _02334_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__a21oi_1
X_08293_ u_rf.reg31_q\[6\] _03289_ _03291_ u_rf.reg11_q\[6\] _03490_ VGND VGND VPWR
+ VPWR _03491_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_621 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07244_ u_rf.reg17_q\[16\] _01630_ _01656_ u_rf.reg10_q\[16\] _02481_ VGND VGND VPWR
+ VPWR _02482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07175_ u_decod.pc_q_o\[15\] _02335_ _01485_ VGND VGND VPWR VPWR _02416_ sky130_fd_sc_hd__o21ai_1
X_06126_ _01359_ _01395_ _01396_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06057_ u_decod.rs2_data_q\[6\] u_decod.rs1_data_q\[6\] VGND VGND VPWR VPWR _01328_
+ sky130_fd_sc_hd__nor2_1
Xfanout301 net310 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_93_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout312 net318 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_4
Xfanout323 net327 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_4
Xfanout356 net358 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_2
Xfanout345 net348 VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__buf_2
XFILLER_0_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout334 net374 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_4
Xfanout367 net373 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_2
X_09816_ u_rf.reg6_q\[8\] _04444_ _04684_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__mux2_1
X_09747_ u_rf.reg5_q\[8\] _04444_ _04647_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__mux2_1
X_06959_ u_rf.reg5_q\[11\] _01568_ _01670_ u_rf.reg27_q\[11\] VGND VGND VPWR VPWR
+ _02207_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_124_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_649 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09678_ u_rf.reg4_q\[9\] _04446_ _04608_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _03805_ _03807_ _03809_ _03811_ VGND VGND VPWR VPWR _03812_ sky130_fd_sc_hd__or4_1
X_11640_ net344 VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11571_ _04568_ _04936_ _05114_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__or3_4
XFILLER_0_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10522_ _05099_ VGND VGND VPWR VPWR _00499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10453_ _04761_ u_rf.reg14_q\[19\] _05053_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10384_ _05026_ VGND VGND VPWR VPWR _00434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12123_ clknet_leaf_10_clk _00160_ net224 VGND VGND VPWR VPWR u_rf.reg5_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_12054_ clknet_leaf_95_clk net437 net333 VGND VGND VPWR VPWR u_decod.rf_ff_rd_adr_q_i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_144_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11005_ u_rf.reg22_q\[21\] _04983_ _05355_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12956_ clknet_leaf_127_clk _00993_ net238 VGND VGND VPWR VPWR u_rf.reg31_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_73_clk _00924_ net359 VGND VGND VPWR VPWR u_rf.reg28_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_11907_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[28\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ clknet_leaf_128_clk _00065_ net236 VGND VGND VPWR VPWR u_rf.reg0_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
X_11769_ clknet_leaf_66_clk _00061_ net355 VGND VGND VPWR VPWR u_rf.reg1_q\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_573 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08980_ _04129_ _04130_ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_58_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07931_ _02621_ _03134_ _03138_ _03139_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07862_ u_rf.reg12_q\[29\] _01610_ _02697_ u_rf.reg4_q\[29\] VGND VGND VPWR VPWR
+ _03074_ sky130_fd_sc_hd__a22o_1
X_09601_ u_rf.reg3_q\[5\] _04438_ _04571_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__mux2_1
X_06813_ u_rf.reg25_q\[8\] _01574_ _01620_ u_rf.reg24_q\[8\] _02066_ VGND VGND VPWR
+ VPWR _02067_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07793_ _02961_ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09532_ _04539_ VGND VGND VPWR VPWR _00069_ sky130_fd_sc_hd__clkbuf_1
X_06744_ _01444_ _02000_ _01497_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09463_ _04502_ VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__clkbuf_1
X_06675_ u_rf.reg13_q\[5\] _01596_ _01626_ u_rf.reg29_q\[5\] VGND VGND VPWR VPWR _01935_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09394_ u_decod.rf_ff_res_data_i\[14\] VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__buf_2
X_08414_ net448 _03565_ _03606_ _03586_ VGND VGND VPWR VPWR u_decod.rs1_data\[11\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_630 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08345_ _03531_ _03540_ _03337_ VGND VGND VPWR VPWR _03541_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_31_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08276_ _03468_ _03470_ _03472_ _03474_ VGND VGND VPWR VPWR _03475_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07227_ u_decod.dec0.instr_i\[16\] _01208_ _02256_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07158_ _01289_ _01447_ _01685_ _02136_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06109_ u_decod.rs1_data_q\[17\] VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07089_ _01437_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_clk clknet_4_10_0_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_126_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12810_ clknet_leaf_27_clk _00847_ net259 VGND VGND VPWR VPWR u_rf.reg26_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ clknet_leaf_121_clk _00778_ net247 VGND VGND VPWR VPWR u_rf.reg24_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12672_ clknet_leaf_119_clk _00709_ net249 VGND VGND VPWR VPWR u_rf.reg22_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11623_ _04772_ u_rf.reg31_q\[24\] _05679_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_721 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11554_ _05647_ VGND VGND VPWR VPWR _00983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11485_ _04770_ u_rf.reg29_q\[23\] _05607_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _04745_ u_rf.reg15_q\[11\] _05089_ VGND VGND VPWR VPWR _05091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_688 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10436_ _05054_ VGND VGND VPWR VPWR _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10367_ _04742_ u_rf.reg13_q\[10\] _05017_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12106_ clknet_leaf_30_clk _00143_ net261 VGND VGND VPWR VPWR u_rf.reg4_q\[15\] sky130_fd_sc_hd__dfrtp_1
X_10298_ u_decod.rf_ff_res_data_i\[17\] VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_287 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_89_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
X_12037_ clknet_leaf_96_clk u_decod.exe_ff_res_data_i\[17\] net331 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12939_ clknet_leaf_136_clk _00976_ net205 VGND VGND VPWR VPWR u_rf.reg30_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_146_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06460_ u_rf.reg25_q\[1\] _01576_ _01630_ u_rf.reg17_q\[1\] _01727_ VGND VGND VPWR
+ VPWR _01728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_157_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
X_08130_ u_rf.reg28_q\[0\] _03331_ _03333_ u_rf.reg2_q\[0\] VGND VGND VPWR VPWR _03334_
+ sky130_fd_sc_hd__a22o_1
X_06391_ u_rf.reg4_q\[0\] _01650_ _01654_ u_rf.reg22_q\[0\] _01660_ VGND VGND VPWR
+ VPWR _01661_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08061_ _03264_ VGND VGND VPWR VPWR _03265_ sky130_fd_sc_hd__buf_8
XFILLER_0_114_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07012_ u_rf.reg25_q\[12\] _01575_ _01624_ u_rf.reg28_q\[12\] VGND VGND VPWR VPWR
+ _02258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08963_ _04101_ _04116_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07914_ _03114_ _03123_ _02359_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__o21a_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08894_ _04050_ net387 _04049_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07845_ _01260_ _03047_ _03055_ _03057_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__a211o_1
X_07776_ _02982_ _02991_ _02359_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_104_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09515_ _04529_ VGND VGND VPWR VPWR _00062_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06727_ u_rf.reg30_q\[6\] _01579_ _01608_ u_rf.reg12_q\[6\] _01984_ VGND VGND VPWR
+ VPWR _01985_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_121_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ u_decod.rf_ff_res_data_i\[31\] VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__buf_2
XFILLER_0_78_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06658_ _01764_ _01917_ _01918_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__or3b_1
XFILLER_0_74_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06589_ _01772_ u_decod.exe_ff_res_data_i\[3\] _01832_ _01852_ VGND VGND VPWR VPWR
+ _01853_ sky130_fd_sc_hd__a211o_1
X_09377_ _04445_ VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08328_ u_rf.reg18_q\[8\] _03262_ _03263_ u_rf.reg23_q\[8\] _03523_ VGND VGND VPWR
+ VPWR _03524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08259_ u_rf.reg12_q\[5\] _03241_ _03202_ u_rf.reg10_q\[5\] VGND VGND VPWR VPWR _03458_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11270_ u_rf.reg26_q\[18\] u_decod.rf_ff_res_data_i\[18\] _05488_ VGND VGND VPWR
+ VPWR _05497_ sky130_fd_sc_hd__mux2_1
X_10221_ _04924_ VGND VGND VPWR VPWR _00373_ sky130_fd_sc_hd__clkbuf_1
X_10152_ _04887_ VGND VGND VPWR VPWR _00341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_440 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10083_ u_rf.reg9_q\[21\] _04472_ _04849_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12724_ clknet_leaf_24_clk _00761_ net267 VGND VGND VPWR VPWR u_rf.reg23_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10985_ _05346_ VGND VGND VPWR VPWR _00715_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ clknet_leaf_37_clk _00692_ net272 VGND VGND VPWR VPWR u_rf.reg21_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12586_ clknet_leaf_29_clk _00623_ net259 VGND VGND VPWR VPWR u_rf.reg19_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11606_ _04755_ u_rf.reg31_q\[16\] _05668_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11537_ _05638_ VGND VGND VPWR VPWR _00975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_705 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11468_ _04753_ u_rf.reg29_q\[15\] _05596_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11399_ _05565_ VGND VGND VPWR VPWR _00910_ sky130_fd_sc_hd__clkbuf_1
X_10419_ _05045_ VGND VGND VPWR VPWR _00450_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
X_05960_ _01088_ VGND VGND VPWR VPWR _01239_ sky130_fd_sc_hd__inv_2
X_05891_ _01099_ _01183_ _01184_ _01185_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07630_ u_rf.reg7_q\[24\] _01562_ _01780_ u_rf.reg29_q\[24\] _02851_ VGND VGND VPWR
+ VPWR _02852_ sky130_fd_sc_hd__a221o_1
X_07561_ _02579_ _02785_ _01464_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_736 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06512_ u_rf.reg31_q\[2\] _01777_ _01650_ u_rf.reg4_q\[2\] VGND VGND VPWR VPWR _01778_
+ sky130_fd_sc_hd__a22o_1
X_09300_ u_decod.instr_unit_q\[3\] VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_152_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07492_ _02718_ _02719_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[21\] sky130_fd_sc_hd__xor2_1
XFILLER_0_146_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09231_ _04342_ _04343_ _04340_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__o21a_1
XFILLER_0_119_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_326 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06443_ _01693_ _01701_ _01711_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__or3_1
X_09162_ _04078_ _04274_ _04275_ _04289_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[14\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_84_791 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06374_ _01643_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__buf_8
XFILLER_0_145_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08113_ u_rf.reg1_q\[0\] _03311_ _03313_ u_rf.reg14_q\[0\] _03316_ VGND VGND VPWR
+ VPWR _03317_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09093_ _04228_ _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08044_ u_rf.reg16_q\[31\] _03248_ _03249_ u_rf.reg5_q\[31\] VGND VGND VPWR VPWR
+ _03250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09995_ u_rf.reg8_q\[12\] _04453_ _04801_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__mux2_1
X_08946_ _01376_ u_decod.branch_imm_q_o\[19\] VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_4_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ u_decod.rs1_data_q\[9\] u_decod.branch_imm_q_o\[9\] VGND VGND VPWR VPWR _04043_
+ sky130_fd_sc_hd__nor2_1
X_07828_ _02994_ _02996_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07759_ u_rf.reg13_q\[27\] _02376_ _01787_ u_rf.reg18_q\[27\] _02974_ VGND VGND VPWR
+ VPWR _02975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10770_ u_rf.reg19_q\[7\] _04953_ _05224_ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__mux2_1
X_09429_ u_rf.reg2_q\[25\] _04480_ _04470_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12440_ clknet_leaf_67_clk _00477_ net349 VGND VGND VPWR VPWR u_rf.reg14_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12371_ clknet_leaf_69_clk _00408_ net350 VGND VGND VPWR VPWR u_rf.reg12_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_134_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11322_ _04742_ u_rf.reg27_q\[10\] _05524_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__mux2_1
X_11253_ _05476_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__buf_6
X_10204_ _04915_ VGND VGND VPWR VPWR _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11184_ _05451_ VGND VGND VPWR VPWR _00809_ sky130_fd_sc_hd__clkbuf_1
X_10135_ _04878_ VGND VGND VPWR VPWR _00333_ sky130_fd_sc_hd__clkbuf_1
X_10066_ u_rf.reg9_q\[13\] _04455_ _04838_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_50_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10968_ _05337_ VGND VGND VPWR VPWR _00707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12707_ clknet_leaf_106_clk _00744_ net319 VGND VGND VPWR VPWR u_rf.reg23_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10899_ u_rf.reg21_q\[3\] _04945_ _05297_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__mux2_1
X_12638_ clknet_leaf_123_clk _00675_ net232 VGND VGND VPWR VPWR u_rf.reg21_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12569_ clknet_leaf_64_clk _00606_ net341 VGND VGND VPWR VPWR u_rf.reg18_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06090_ _01359_ _01360_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08800_ u_decod.rf_ff_res_data_i\[29\] _03382_ _03974_ _03404_ VGND VGND VPWR VPWR
+ _03975_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09780_ _04673_ VGND VGND VPWR VPWR _00183_ sky130_fd_sc_hd__clkbuf_1
X_06992_ _02038_ _02238_ _01451_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08731_ u_rf.reg16_q\[26\] _03450_ _03515_ u_rf.reg5_q\[26\] VGND VGND VPWR VPWR
+ _03909_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_0_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_05943_ _01202_ u_decod.dec0.is_shift _01224_ VGND VGND VPWR VPWR u_decod.dec0.is_arithm
+ sky130_fd_sc_hd__o21bai_1
X_08662_ u_rf.reg30_q\[23\] _03281_ _03283_ u_rf.reg10_q\[23\] _03842_ VGND VGND VPWR
+ VPWR _03843_ sky130_fd_sc_hd__a221o_1
X_05874_ _01171_ _01144_ _01172_ VGND VGND VPWR VPWR _01173_ sky130_fd_sc_hd__and3b_1
X_07613_ _02779_ _02835_ _01480_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__mux2_1
X_08593_ u_rf.reg8_q\[20\] _03271_ _03273_ u_rf.reg29_q\[20\] _03776_ VGND VGND VPWR
+ VPWR _03777_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07544_ _02768_ _02769_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[22\] sky130_fd_sc_hd__nor2_1
XFILLER_0_48_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07475_ u_rf.reg11_q\[21\] _01584_ _01667_ u_rf.reg8_q\[21\] _02702_ VGND VGND VPWR
+ VPWR _02703_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09214_ _04123_ _04206_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06426_ _01314_ _01316_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_249 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09145_ _04206_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06357_ _01626_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_116_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09076_ u_decod.pc_q_o\[3\] u_decod.branch_imm_q_o\[3\] VGND VGND VPWR VPWR _04215_
+ sky130_fd_sc_hd__nor2_1
X_06288_ _01520_ _01552_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__nor2_2
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08027_ u_rf.reg1_q\[31\] _03231_ _03232_ u_rf.reg14_q\[31\] VGND VGND VPWR VPWR
+ _03233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09978_ u_rf.reg8_q\[4\] _04436_ _04790_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__mux2_1
X_08929_ _01292_ u_decod.branch_imm_q_o\[14\] _04087_ _04080_ VGND VGND VPWR VPWR
+ _04088_ sky130_fd_sc_hd__a31o_1
X_11940_ clknet_leaf_74_clk u_decod.rs1_data\[28\] net357 VGND VGND VPWR VPWR u_decod.rs1_data_q\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ clknet_leaf_102_clk u_decod.dec0.operation_o\[2\] net337 VGND VGND VPWR VPWR
+ u_decod.instr_operation_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_10822_ _04606_ _05114_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10753_ _05222_ VGND VGND VPWR VPWR _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10684_ u_rf.reg17_q\[31\] _05003_ _05151_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_457 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12423_ clknet_leaf_3_clk _00460_ net213 VGND VGND VPWR VPWR u_rf.reg14_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_660 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12354_ clknet_leaf_130_clk _00391_ net229 VGND VGND VPWR VPWR u_rf.reg12_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11305_ _04726_ u_rf.reg27_q\[2\] _05513_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12285_ clknet_leaf_14_clk _00322_ net246 VGND VGND VPWR VPWR u_rf.reg10_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11236_ _05479_ VGND VGND VPWR VPWR _00833_ sky130_fd_sc_hd__clkbuf_1
X_11167_ u_rf.reg25_q\[1\] _04941_ _05441_ VGND VGND VPWR VPWR _05443_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10118_ _04869_ VGND VGND VPWR VPWR _00325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11098_ _05406_ VGND VGND VPWR VPWR _00768_ sky130_fd_sc_hd__clkbuf_1
X_10049_ u_rf.reg9_q\[5\] _04438_ _04827_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_717 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07260_ _02189_ _02495_ _02496_ _01441_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07191_ u_rf.reg29_q\[15\] _01628_ _01653_ u_rf.reg22_q\[15\] VGND VGND VPWR VPWR
+ _02431_ sky130_fd_sc_hd__a22o_1
X_06211_ _01452_ _01459_ _01465_ _01473_ _01477_ _01481_ VGND VGND VPWR VPWR _01482_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06142_ _01284_ _01412_ _01281_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06073_ u_decod.rs2_data_q\[10\] _01302_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_343 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09901_ _04742_ u_rf.reg7_q\[10\] _04743_ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09832_ _04701_ VGND VGND VPWR VPWR _00207_ sky130_fd_sc_hd__clkbuf_1
X_09763_ _04664_ VGND VGND VPWR VPWR _00175_ sky130_fd_sc_hd__clkbuf_1
X_08714_ _03886_ _03888_ _03890_ _03892_ VGND VGND VPWR VPWR _03893_ sky130_fd_sc_hd__or4_1
X_06975_ _02213_ _02222_ _01679_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__o21a_2
Xrebuffer21 net396 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 _01124_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
X_09694_ _04626_ VGND VGND VPWR VPWR _00144_ sky130_fd_sc_hd__clkbuf_1
X_05926_ _01214_ VGND VGND VPWR VPWR u_decod.dec0.rd_o\[0\] sky130_fd_sc_hd__clkbuf_1
Xrebuffer32 _04164_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
X_05857_ u_decod.pc0_q_i\[17\] u_decod.pc0_q_i\[18\] _01150_ u_decod.pc0_q_i\[19\]
+ VGND VGND VPWR VPWR _01160_ sky130_fd_sc_hd__a31o_1
X_08645_ u_rf.reg6_q\[22\] _03387_ _03344_ u_rf.reg26_q\[22\] _03826_ VGND VGND VPWR
+ VPWR _03827_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_820 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08576_ u_rf.reg26_q\[19\] _03343_ _03285_ u_rf.reg21_q\[19\] VGND VGND VPWR VPWR
+ _03761_ sky130_fd_sc_hd__a22o_1
X_07527_ _02746_ _02748_ _02750_ _02752_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__or4_1
X_05788_ net480 _01105_ _01101_ net87 _01107_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__a221o_1
XFILLER_0_37_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07458_ _02631_ _02686_ _02189_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_295 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07389_ _02619_ net45 VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06409_ _01678_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_400 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09128_ _04253_ _04248_ _04250_ _04251_ _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__o311a_1
XFILLER_0_17_485 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_855 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09059_ _01066_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12070_ clknet_leaf_140_clk _00107_ net202 VGND VGND VPWR VPWR u_rf.reg3_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11021_ u_rf.reg22_q\[29\] _04999_ _05355_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12972_ clknet_leaf_14_clk _01009_ net246 VGND VGND VPWR VPWR u_rf.reg31_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11923_ clknet_leaf_87_clk u_decod.rs1_data\[11\] net362 VGND VGND VPWR VPWR u_decod.rs1_data_q\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_142_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ clknet_leaf_14_clk _00081_ net244 VGND VGND VPWR VPWR u_rf.reg0_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_10805_ _05250_ VGND VGND VPWR VPWR _00631_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11785_ clknet_leaf_84_clk net137 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_694 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10736_ u_rf.reg18_q\[23\] _04987_ _05210_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_322 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10667_ _05177_ VGND VGND VPWR VPWR _00566_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12406_ clknet_leaf_49_clk _00443_ net306 VGND VGND VPWR VPWR u_rf.reg13_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10598_ u_rf.reg16_q\[22\] _04985_ _05138_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net119 VGND VGND VPWR VPWR adr_o[26] sky130_fd_sc_hd__buf_4
Xoutput108 net108 VGND VGND VPWR VPWR adr_o[16] sky130_fd_sc_hd__buf_4
X_12337_ clknet_leaf_22_clk _00374_ net285 VGND VGND VPWR VPWR u_rf.reg11_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_81_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ clknet_leaf_14_clk _00305_ net244 VGND VGND VPWR VPWR u_rf.reg9_q\[17\] sky130_fd_sc_hd__dfrtp_1
X_11219_ u_rf.reg25_q\[26\] _04993_ _05463_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__mux2_1
X_12199_ clknet_leaf_3_clk _00236_ net213 VGND VGND VPWR VPWR u_rf.reg7_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06760_ u_rf.reg16_q\[7\] _01563_ _01651_ u_rf.reg22_q\[7\] VGND VGND VPWR VPWR _02016_
+ sky130_fd_sc_hd__a22o_1
X_06691_ u_decod.rs1_data_q\[21\] _01446_ _01753_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_90_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08430_ u_rf.reg28_q\[12\] _03331_ _03557_ u_rf.reg2_q\[12\] VGND VGND VPWR VPWR
+ _03622_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_503 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08361_ _03330_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__buf_8
XFILLER_0_129_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08292_ u_rf.reg9_q\[6\] _03212_ _03213_ u_rf.reg20_q\[6\] VGND VGND VPWR VPWR _03490_
+ sky130_fd_sc_hd__a22o_1
X_07312_ _01403_ _01429_ _02539_ _02545_ _02546_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_144_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07243_ u_rf.reg29_q\[16\] _01627_ _01652_ u_rf.reg22_q\[16\] VGND VGND VPWR VPWR
+ _02481_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_720 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07174_ _01746_ _02402_ _02409_ _02414_ VGND VGND VPWR VPWR _02415_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06125_ u_decod.rs2_data_q\[21\] _01358_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06056_ _01325_ _01326_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__nor2_1
Xfanout302 net305 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout313 net318 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_4
Xfanout357 net358 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
Xfanout346 net348 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_4
Xfanout324 net327 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_4
X_09815_ _04692_ VGND VGND VPWR VPWR _00199_ sky130_fd_sc_hd__clkbuf_1
Xfanout335 net336 VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_4
Xfanout368 net373 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_129_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09746_ _04655_ VGND VGND VPWR VPWR _00167_ sky130_fd_sc_hd__clkbuf_1
X_06958_ u_rf.reg31_q\[11\] _01616_ _01639_ u_rf.reg21_q\[11\] _02205_ VGND VGND VPWR
+ VPWR _02206_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09677_ _04617_ VGND VGND VPWR VPWR _00136_ sky130_fd_sc_hd__clkbuf_1
X_05909_ u_decod.dec0.instr_i\[0\] _01074_ VGND VGND VPWR VPWR _01199_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_124_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ u_rf.reg27_q\[21\] _03319_ _03321_ u_rf.reg19_q\[21\] _03810_ VGND VGND VPWR
+ VPWR _03811_ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06889_ _02102_ _02139_ _01422_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_38_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08559_ u_rf.reg15_q\[18\] _03237_ _03302_ u_rf.reg24_q\[18\] VGND VGND VPWR VPWR
+ _03745_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11570_ _05655_ VGND VGND VPWR VPWR _00991_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ _04761_ u_rf.reg15_q\[19\] _05089_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_138_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10452_ _05062_ VGND VGND VPWR VPWR _00466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10383_ _04759_ u_rf.reg13_q\[18\] _05017_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12122_ clknet_leaf_59_clk _00159_ net289 VGND VGND VPWR VPWR u_rf.reg4_q\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12053_ clknet_leaf_95_clk net447 net325 VGND VGND VPWR VPWR u_decod.rf_ff_rd_adr_q_i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_11004_ _05356_ VGND VGND VPWR VPWR _00724_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ clknet_leaf_122_clk _00992_ net242 VGND VGND VPWR VPWR u_rf.reg31_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11906_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[27\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ clknet_leaf_73_clk _00923_ net359 VGND VGND VPWR VPWR u_rf.reg28_q\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_138 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11837_ clknet_leaf_13_clk _00064_ net244 VGND VGND VPWR VPWR u_rf.reg0_q\[0\] sky130_fd_sc_hd__dfrtp_1
X_11768_ clknet_leaf_71_clk _00060_ net358 VGND VGND VPWR VPWR u_rf.reg1_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10719_ u_rf.reg18_q\[15\] _04970_ _05199_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11699_ _05724_ VGND VGND VPWR VPWR _01051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_788 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_585 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer1 u_decod.rs1_data_q\[1\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07930_ _02789_ _03099_ _01507_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_58_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07861_ u_rf.reg15_q\[29\] _02371_ _02379_ u_rf.reg17_q\[29\] _03072_ VGND VGND VPWR
+ VPWR _03073_ sky130_fd_sc_hd__a221o_1
X_07792_ _02619_ net53 _02618_ VGND VGND VPWR VPWR _03007_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09600_ _04576_ VGND VGND VPWR VPWR _00100_ sky130_fd_sc_hd__clkbuf_1
X_06812_ u_rf.reg26_q\[8\] _01640_ _01643_ u_rf.reg20_q\[8\] VGND VGND VPWR VPWR _02066_
+ sky130_fd_sc_hd__a22o_1
X_09531_ u_rf.reg0_q\[5\] _04438_ _04533_ VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__mux2_1
X_06743_ u_decod.rs1_data_q\[7\] _01702_ _01703_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09462_ u_rf.reg1_q\[5\] _04438_ _04496_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__mux2_1
X_06674_ u_rf.reg16_q\[5\] _01564_ _01615_ u_rf.reg31_q\[5\] _01933_ VGND VGND VPWR
+ VPWR _01934_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09393_ _04456_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__clkbuf_1
X_08413_ u_decod.exe_ff_res_data_i\[11\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[11\]
+ _03605_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__a221o_2
XFILLER_0_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08344_ _03533_ _03535_ _03537_ _03539_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08275_ u_rf.reg18_q\[5\] _03262_ _03366_ u_rf.reg19_q\[5\] _03473_ VGND VGND VPWR
+ VPWR _03474_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07226_ _01437_ _02442_ _02443_ _02464_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[16\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07157_ _02397_ _01352_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06108_ _01377_ _01378_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07088_ _01295_ _01299_ _01351_ _01355_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__o31ai_2
X_06039_ u_decod.rs2_data_q\[5\] u_decod.rs1_data_q\[5\] VGND VGND VPWR VPWR _01310_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ _04643_ _04644_ _04645_ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__and3_4
XFILLER_0_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ clknet_leaf_112_clk _00777_ net317 VGND VGND VPWR VPWR u_rf.reg24_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12671_ clknet_leaf_137_clk _00708_ net205 VGND VGND VPWR VPWR u_rf.reg22_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11622_ _05683_ VGND VGND VPWR VPWR _01015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_146_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _04770_ u_rf.reg30_q\[23\] _05643_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11484_ _05610_ VGND VGND VPWR VPWR _00950_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10504_ _05090_ VGND VGND VPWR VPWR _00490_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_555 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10435_ _04742_ u_rf.reg14_q\[10\] _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_572 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12105_ clknet_leaf_23_clk _00142_ net284 VGND VGND VPWR VPWR u_rf.reg4_q\[14\] sky130_fd_sc_hd__dfrtp_1
X_10366_ _05005_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__buf_6
XPHY_EDGE_ROW_155_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10297_ _04973_ VGND VGND VPWR VPWR _00400_ sky130_fd_sc_hd__clkbuf_1
X_12036_ clknet_leaf_95_clk u_decod.exe_ff_res_data_i\[16\] net331 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_88_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12938_ clknet_leaf_30_clk _00975_ net262 VGND VGND VPWR VPWR u_rf.reg30_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_157_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12869_ clknet_leaf_121_clk _00906_ net249 VGND VGND VPWR VPWR u_rf.reg28_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06390_ u_rf.reg10_q\[0\] _01656_ _01659_ u_rf.reg14_q\[0\] VGND VGND VPWR VPWR _01660_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08060_ _03224_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__buf_6
XFILLER_0_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07011_ u_decod.dec0.funct3\[0\] _01208_ _02256_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__a21o_2
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ _04114_ _04115_ VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_90_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07913_ _03116_ _03118_ _03120_ _03122_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__or4_1
X_08893_ _04055_ _04056_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__nor2_1
X_07844_ u_decod.pc_q_o\[29\] _02999_ _03056_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07775_ _02984_ _02986_ _02988_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09514_ u_rf.reg1_q\[30\] _04490_ _04495_ VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_918 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06726_ u_rf.reg24_q\[6\] _01621_ _01624_ u_rf.reg28_q\[6\] VGND VGND VPWR VPWR _01984_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _04491_ VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06657_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] u_decod.pc_q_o\[4\] u_decod.pc_q_o\[5\]
+ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06588_ _01680_ _01851_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__and2_1
X_09376_ u_rf.reg2_q\[8\] _04444_ _04428_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__mux2_1
X_08327_ u_rf.reg4_q\[8\] _03265_ _03267_ u_rf.reg17_q\[8\] VGND VGND VPWR VPWR _03523_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08258_ net386 _03259_ _03457_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[4\]
+ sky130_fd_sc_hd__a22o_1
X_07209_ _02446_ _02447_ _01057_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10220_ _04766_ u_rf.reg11_q\[21\] _04922_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__mux2_1
X_08189_ u_rf.reg16_q\[2\] _03322_ _03324_ u_rf.reg5_q\[2\] VGND VGND VPWR VPWR _03391_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10151_ u_rf.reg10_q\[21\] _04472_ _04885_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10082_ _04850_ VGND VGND VPWR VPWR _00308_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_531 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10984_ u_rf.reg22_q\[11\] _04962_ _05344_ VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__mux2_1
X_12723_ clknet_leaf_52_clk _00760_ net351 VGND VGND VPWR VPWR u_rf.reg23_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ clknet_leaf_7_clk _00691_ net219 VGND VGND VPWR VPWR u_rf.reg21_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12585_ clknet_leaf_25_clk _00622_ net280 VGND VGND VPWR VPWR u_rf.reg19_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_11605_ _05674_ VGND VGND VPWR VPWR _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11536_ _04753_ u_rf.reg30_q\[15\] _05632_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_291 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_152_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11467_ _05601_ VGND VGND VPWR VPWR _00942_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11398_ net525 u_decod.rf_ff_res_data_i\[14\] _05560_ VGND VGND VPWR VPWR _05565_
+ sky130_fd_sc_hd__mux2_1
X_10418_ _04726_ u_rf.reg14_q\[2\] _05042_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _05008_ VGND VGND VPWR VPWR _00417_ sky130_fd_sc_hd__clkbuf_1
X_12019_ clknet_leaf_97_clk net476 net332 VGND VGND VPWR VPWR u_exe.flush_v_dly1_q
+ sky130_fd_sc_hd__dfrtp_1
X_05890_ u_exe.pc_data_q\[27\] _01118_ _01100_ net84 VGND VGND VPWR VPWR _01185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07560_ _01467_ _02404_ _01498_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__o21a_1
X_06511_ _01616_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09230_ _04345_ _04346_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__nand2_1
X_07491_ _01897_ _02671_ _02673_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_625 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06442_ _01505_ _01708_ _01710_ _01058_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09161_ _04287_ _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_483 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06373_ _01538_ _01514_ _01551_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__and3_2
X_09092_ _04223_ _04224_ _04221_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__o21a_1
X_08112_ u_rf.reg7_q\[0\] _03314_ _03315_ u_rf.reg25_q\[0\] VGND VGND VPWR VPWR _03316_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_133 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08043_ _03170_ _03204_ _03205_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__and3_4
XFILLER_0_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_238 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09994_ _04803_ VGND VGND VPWR VPWR _00267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08945_ _02621_ VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_4_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08876_ _02621_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07827_ _02357_ u_decod.exe_ff_res_data_i\[28\] _03040_ VGND VGND VPWR VPWR _03041_
+ sky130_fd_sc_hd__a21o_1
X_07758_ u_rf.reg27_q\[27\] _02386_ _01776_ u_rf.reg2_q\[27\] VGND VGND VPWR VPWR
+ _02974_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06709_ _01765_ _01948_ _01954_ _01967_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__o211a_1
X_07689_ u_decod.pc_q_o\[26\] _02868_ VGND VGND VPWR VPWR _02908_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ u_decod.rf_ff_res_data_i\[25\] VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_23_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09359_ _04433_ VGND VGND VPWR VPWR _00002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ clknet_leaf_41_clk _00407_ net277 VGND VGND VPWR VPWR u_rf.reg12_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11321_ _05512_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_134_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11252_ _05487_ VGND VGND VPWR VPWR _00841_ sky130_fd_sc_hd__clkbuf_1
X_10203_ _04749_ u_rf.reg11_q\[13\] _04911_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__mux2_1
X_11183_ u_rf.reg25_q\[9\] _04957_ _05441_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10134_ u_rf.reg10_q\[13\] _04455_ _04874_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__mux2_1
X_10065_ _04841_ VGND VGND VPWR VPWR _00300_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10967_ u_rf.reg22_q\[3\] _04945_ _05333_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10898_ _05300_ VGND VGND VPWR VPWR _00674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12706_ clknet_leaf_130_clk _00743_ net229 VGND VGND VPWR VPWR u_rf.reg23_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12637_ clknet_leaf_16_clk _00674_ net250 VGND VGND VPWR VPWR u_rf.reg21_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12568_ clknet_leaf_68_clk _00605_ net351 VGND VGND VPWR VPWR u_rf.reg18_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12499_ clknet_leaf_68_clk _00536_ net350 VGND VGND VPWR VPWR u_rf.reg16_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11519_ _04736_ u_rf.reg30_q\[7\] _05621_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06991_ _02236_ _02237_ _01455_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08730_ u_rf.reg7_q\[26\] _03369_ _03370_ u_rf.reg25_q\[26\] _03907_ VGND VGND VPWR
+ VPWR _03908_ sky130_fd_sc_hd__a221o_1
X_05942_ _01206_ VGND VGND VPWR VPWR _01224_ sky130_fd_sc_hd__clkbuf_4
X_08661_ u_rf.reg26_q\[23\] _03284_ _03286_ u_rf.reg21_q\[23\] VGND VGND VPWR VPWR
+ _03842_ sky130_fd_sc_hd__a22o_1
X_05873_ u_decod.pc0_q_i\[23\] _01168_ VGND VGND VPWR VPWR _01172_ sky130_fd_sc_hd__or2_1
X_07612_ _02733_ _02834_ _01476_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__mux2_1
X_08592_ u_rf.reg22_q\[20\] _03409_ _03277_ u_rf.reg3_q\[20\] VGND VGND VPWR VPWR
+ _03776_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07543_ _02765_ _02767_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07474_ u_rf.reg6_q\[21\] _01556_ _01653_ u_rf.reg22_q\[21\] VGND VGND VPWR VPWR
+ _02702_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09213_ _04330_ _04332_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06425_ _01314_ _01316_ VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09144_ _04066_ _04207_ _04208_ _04273_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[12\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_101_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06356_ _01572_ _01566_ _01577_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__and3_2
XFILLER_0_126_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09075_ _04198_ _04202_ _04203_ _04211_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__o211a_1
X_06287_ _01556_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_8
X_08026_ _03170_ _03198_ _03199_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__and3_4
XFILLER_0_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09977_ _04794_ VGND VGND VPWR VPWR _00259_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_110_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08928_ _01289_ u_decod.branch_imm_q_o\[15\] VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08859_ _04014_ _04016_ _04020_ _04027_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_28_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11870_ clknet_leaf_103_clk u_decod.dec0.operation_o\[1\] net336 VGND VGND VPWR VPWR
+ u_decod.instr_operation_q\[1\] sky130_fd_sc_hd__dfrtp_4
X_10821_ _05258_ VGND VGND VPWR VPWR _00639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10752_ u_rf.reg18_q\[31\] _05003_ _05187_ VGND VGND VPWR VPWR _05222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10683_ _05185_ VGND VGND VPWR VPWR _00574_ sky130_fd_sc_hd__clkbuf_1
X_12422_ clknet_leaf_140_clk _00459_ net203 VGND VGND VPWR VPWR u_rf.reg14_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_801 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12353_ clknet_leaf_119_clk _00390_ net251 VGND VGND VPWR VPWR u_rf.reg12_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11304_ _05515_ VGND VGND VPWR VPWR _00865_ sky130_fd_sc_hd__clkbuf_1
X_12284_ clknet_leaf_127_clk _00321_ net237 VGND VGND VPWR VPWR u_rf.reg10_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_309 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11235_ u_rf.reg26_q\[1\] net496 _05477_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ _05442_ VGND VGND VPWR VPWR _00800_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11097_ u_rf.reg24_q\[0\] _04935_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__mux2_1
X_10117_ u_rf.reg10_q\[5\] _04438_ _04863_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10048_ _04832_ VGND VGND VPWR VPWR _00292_ sky130_fd_sc_hd__clkbuf_1
Xhold90 u_decod.pc0_q_i\[26\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11999_ clknet_leaf_82_clk u_exe.bu_pc_res\[12\] net364 VGND VGND VPWR VPWR u_exe.pc_data_q\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06210_ _01480_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_303 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07190_ u_rf.reg11_q\[15\] _01584_ _02376_ u_rf.reg13_q\[15\] _02429_ VGND VGND VPWR
+ VPWR _02430_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06141_ _01409_ _01411_ _01282_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__o21a_1
XFILLER_0_54_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06072_ u_decod.rs2_data_q\[10\] u_decod.rs1_data_q\[10\] VGND VGND VPWR VPWR _01343_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_467 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09900_ _04721_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ u_rf.reg6_q\[15\] _04459_ _04695_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09762_ u_rf.reg5_q\[15\] _04459_ _04658_ VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__mux2_1
X_06974_ _02215_ _02217_ _02219_ _02221_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__or4_1
X_08713_ u_rf.reg16_q\[25\] _03323_ _03325_ u_rf.reg5_q\[25\] _03891_ VGND VGND VPWR
+ VPWR _03892_ sky130_fd_sc_hd__a221o_1
X_05925_ u_decod.dec0.instr_i\[7\] u_decod.dec0.rd_v VGND VGND VPWR VPWR _01214_ sky130_fd_sc_hd__and2_1
Xrebuffer11 net410 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09693_ u_rf.reg4_q\[16\] _04461_ _04619_ VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__mux2_1
X_05856_ u_decod.pc0_q_i\[18\] u_decod.pc0_q_i\[19\] _01153_ VGND VGND VPWR VPWR _01159_
+ sky130_fd_sc_hd__and3_1
Xrebuffer22 net397 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
X_08644_ u_rf.reg18_q\[22\] _03222_ _03223_ u_rf.reg23_q\[22\] VGND VGND VPWR VPWR
+ _03826_ sky130_fd_sc_hd__a22o_1
Xrebuffer33 _04016_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_05787_ net390 _01106_ VGND VGND VPWR VPWR _01107_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08575_ u_rf.reg31_q\[19\] _03504_ _03505_ u_rf.reg11_q\[19\] _03759_ VGND VGND VPWR
+ VPWR _03760_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07526_ u_rf.reg16_q\[22\] _02307_ _02376_ u_rf.reg13_q\[22\] _02751_ VGND VGND VPWR
+ VPWR _02752_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_879 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07457_ _02400_ _02498_ _02584_ _02684_ _01475_ _02685_ VGND VGND VPWR VPWR _02686_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07388_ net100 VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__buf_2
X_06408_ _01547_ _01517_ _01527_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__and3b_2
XFILLER_0_9_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09127_ _04250_ u_decod.branch_imm_q_o\[8\] u_decod.pc_q_o\[8\] VGND VGND VPWR VPWR
+ _04259_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06339_ _01608_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_131_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09058_ _04194_ _02334_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__nor2_2
XFILLER_0_60_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_434 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08009_ u_rf.reg31_q\[31\] _03210_ _03211_ u_rf.reg11_q\[31\] _03214_ VGND VGND VPWR
+ VPWR _03215_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_489 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11020_ _05364_ VGND VGND VPWR VPWR _00732_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ clknet_leaf_136_clk _01008_ net205 VGND VGND VPWR VPWR u_rf.reg31_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11922_ clknet_leaf_96_clk u_decod.rs1_data\[10\] net333 VGND VGND VPWR VPWR u_decod.rs1_data_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_142_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11853_ clknet_leaf_1_clk _00080_ net208 VGND VGND VPWR VPWR u_rf.reg0_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_517 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10804_ u_rf.reg19_q\[23\] _04987_ _05246_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11784_ clknet_leaf_84_clk net136 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10735_ _05213_ VGND VGND VPWR VPWR _00598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_172 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10666_ u_rf.reg17_q\[22\] _04985_ _05174_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12405_ clknet_leaf_46_clk _00442_ net298 VGND VGND VPWR VPWR u_rf.reg13_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10597_ _05140_ VGND VGND VPWR VPWR _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput109 net109 VGND VGND VPWR VPWR adr_o[17] sky130_fd_sc_hd__buf_2
X_12336_ clknet_leaf_43_clk _00373_ net275 VGND VGND VPWR VPWR u_rf.reg11_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12267_ clknet_leaf_135_clk _00304_ net209 VGND VGND VPWR VPWR u_rf.reg9_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11218_ _05469_ VGND VGND VPWR VPWR _00825_ sky130_fd_sc_hd__clkbuf_1
X_12198_ clknet_leaf_140_clk _00235_ net203 VGND VGND VPWR VPWR u_rf.reg7_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11149_ u_rf.reg24_q\[25\] _04991_ _05427_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06690_ u_decod.rs1_data_q\[13\] u_decod.rs1_data_q\[29\] _01702_ VGND VGND VPWR
+ VPWR _01949_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_82_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08360_ u_rf.reg6_q\[9\] _03387_ _03388_ u_rf.reg13_q\[9\] _03554_ VGND VGND VPWR
+ VPWR _03555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07311_ _01387_ _02244_ _01432_ _01385_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_515 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08291_ u_rf.reg30_q\[6\] _03200_ _03282_ u_rf.reg10_q\[6\] _03488_ VGND VGND VPWR
+ VPWR _03489_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07242_ u_rf.reg11_q\[16\] _01583_ _01597_ u_rf.reg13_q\[16\] _02479_ VGND VGND VPWR
+ VPWR _02480_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07173_ _01290_ _01429_ _02410_ _01059_ _02413_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_299 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06124_ u_decod.rs2_data_q\[20\] _01363_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06055_ u_decod.rs2_data_q\[7\] u_decod.rs1_data_q\[7\] VGND VGND VPWR VPWR _01326_
+ sky130_fd_sc_hd__and2_1
Xfanout303 net305 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_111_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout314 net318 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_4
Xfanout347 net348 VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_4
Xfanout325 net327 VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_4
X_09814_ u_rf.reg6_q\[7\] _04442_ _04684_ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__mux2_1
Xfanout336 net337 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_2
Xfanout369 net373 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_4
Xfanout358 net359 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_4
X_09745_ u_rf.reg5_q\[7\] _04442_ _04647_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__mux2_1
X_06957_ u_rf.reg13_q\[11\] _01597_ _01666_ u_rf.reg8_q\[11\] VGND VGND VPWR VPWR
+ _02205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06888_ _02039_ _02138_ _01493_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__mux2_1
X_09676_ u_rf.reg4_q\[8\] _04444_ _04608_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__mux2_1
X_05908_ _01071_ _01197_ VGND VGND VPWR VPWR _01198_ sky130_fd_sc_hd__nor2_1
X_08627_ u_rf.reg16_q\[21\] _03323_ _03325_ u_rf.reg5_q\[21\] VGND VGND VPWR VPWR
+ _03810_ sky130_fd_sc_hd__a22o_1
X_05839_ net460 _01142_ _01132_ net70 _01146_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_38_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08558_ u_rf.reg19_q\[18\] _03320_ _03270_ u_rf.reg8_q\[18\] _03743_ VGND VGND VPWR
+ VPWR _03744_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08489_ u_rf.reg30_q\[15\] _03341_ _03342_ u_rf.reg10_q\[15\] _03677_ VGND VGND VPWR
+ VPWR _03678_ sky130_fd_sc_hd__a221o_1
X_07509_ net133 _02731_ _02735_ _01746_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10520_ _05098_ VGND VGND VPWR VPWR _00498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10451_ _04759_ u_rf.reg14_q\[18\] _05053_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10382_ _05025_ VGND VGND VPWR VPWR _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12121_ clknet_leaf_56_clk _00158_ net291 VGND VGND VPWR VPWR u_rf.reg4_q\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12052_ clknet_leaf_95_clk u_decod.exe_ff_write_v_q_i net333 VGND VGND VPWR VPWR
+ u_decod.rf_write_v_q_i sky130_fd_sc_hd__dfrtp_1
X_11003_ u_rf.reg22_q\[20\] _04980_ _05355_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ clknet_leaf_61_clk _00991_ net340 VGND VGND VPWR VPWR u_rf.reg30_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11905_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[26\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[26\] sky130_fd_sc_hd__dfrtp_1
X_12885_ clknet_leaf_54_clk _00922_ net303 VGND VGND VPWR VPWR u_rf.reg28_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11836_ clknet_leaf_105_clk net25 net321 VGND VGND VPWR VPWR u_decod.dec0.funct7\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_11767_ clknet_leaf_48_clk _00059_ net306 VGND VGND VPWR VPWR u_rf.reg1_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10718_ _05204_ VGND VGND VPWR VPWR _00590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11698_ u_decod.branch_imm_q_o\[27\] _02973_ _05717_ VGND VGND VPWR VPWR _05724_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_597 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10649_ u_rf.reg17_q\[14\] _04968_ _05163_ VGND VGND VPWR VPWR _05168_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer2 net409 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12319_ clknet_leaf_131_clk _00356_ net227 VGND VGND VPWR VPWR u_rf.reg11_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07860_ u_rf.reg1_q\[29\] _02604_ _02367_ u_rf.reg14_q\[29\] VGND VGND VPWR VPWR
+ _03072_ sky130_fd_sc_hd__a22o_1
X_07791_ _01265_ _03001_ _03004_ _03005_ VGND VGND VPWR VPWR _03006_ sky130_fd_sc_hd__a2bb2o_1
X_06811_ u_rf.reg13_q\[8\] _01596_ _01590_ u_rf.reg18_q\[8\] _02064_ VGND VGND VPWR
+ VPWR _02065_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09530_ _04538_ VGND VGND VPWR VPWR _00068_ sky130_fd_sc_hd__clkbuf_1
X_06742_ _01866_ _01957_ _01476_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09461_ _04501_ VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06673_ u_rf.reg12_q\[5\] _01607_ _01637_ u_rf.reg21_q\[5\] VGND VGND VPWR VPWR _01933_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09392_ u_rf.reg2_q\[13\] _04455_ _04449_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08412_ _03595_ _03604_ _03337_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__o21a_2
XFILLER_0_86_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08343_ u_rf.reg7_q\[8\] _03428_ _03429_ u_rf.reg25_q\[8\] _03538_ VGND VGND VPWR
+ VPWR _03539_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08274_ u_rf.reg0_q\[5\] _03174_ _03285_ u_rf.reg21_q\[5\] VGND VGND VPWR VPWR _03473_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07225_ _02448_ _02460_ _02463_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__or3b_1
XFILLER_0_144_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07156_ _01293_ _02331_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07087_ _01355_ _01295_ _01299_ _01351_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__nor4_1
X_06107_ u_decod.rs2_data_q\[19\] _01376_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06038_ u_decod.rs2_data_q\[5\] u_decod.rs1_data_q\[5\] VGND VGND VPWR VPWR _01309_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_126_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07989_ _01535_ u_decod.dec0.instr_i\[18\] _01544_ _03193_ _03194_ VGND VGND VPWR
+ VPWR _03195_ sky130_fd_sc_hd__a2111o_1
X_09728_ _01532_ _01536_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09659_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__buf_6
X_12670_ clknet_leaf_12_clk _00707_ net243 VGND VGND VPWR VPWR u_rf.reg22_q\[3\] sky130_fd_sc_hd__dfrtp_1
X_11621_ _04770_ u_rf.reg31_q\[23\] _05679_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _05646_ VGND VGND VPWR VPWR _00982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_564 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11483_ _04768_ u_rf.reg29_q\[22\] _05607_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__mux2_1
X_10503_ _04742_ u_rf.reg15_q\[10\] _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10434_ _05041_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_21_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10365_ _05016_ VGND VGND VPWR VPWR _00425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12104_ clknet_leaf_19_clk _00141_ net281 VGND VGND VPWR VPWR u_rf.reg4_q\[13\] sky130_fd_sc_hd__dfrtp_1
X_10296_ u_rf.reg12_q\[16\] _04972_ _04960_ VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12035_ clknet_leaf_93_clk u_decod.exe_ff_res_data_i\[15\] net344 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[15\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12937_ clknet_leaf_22_clk _00974_ net284 VGND VGND VPWR VPWR u_rf.reg30_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_779 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12868_ clknet_leaf_112_clk _00905_ net317 VGND VGND VPWR VPWR u_rf.reg28_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11819_ clknet_leaf_105_clk net6 net319 VGND VGND VPWR VPWR u_decod.dec0.funct3\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_157_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_676 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_239 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12799_ clknet_leaf_132_clk _00836_ net228 VGND VGND VPWR VPWR u_rf.reg26_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_372 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07010_ _01226_ _01530_ u_decod.dec0.funct7\[6\] VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__o21a_4
XFILLER_0_113_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08961_ _04108_ _04111_ _04106_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_90_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07912_ u_rf.reg21_q\[30\] _02364_ _02367_ u_rf.reg14_q\[30\] _03121_ VGND VGND VPWR
+ VPWR _03122_ sky130_fd_sc_hd__a221o_1
X_08892_ u_decod.rs1_data_q\[11\] u_decod.branch_imm_q_o\[11\] VGND VGND VPWR VPWR
+ _04056_ sky130_fd_sc_hd__and2_1
X_07843_ u_decod.pc_q_o\[29\] _02999_ _01485_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_108_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07774_ u_rf.reg25_q\[27\] _01783_ _01784_ u_rf.reg24_q\[27\] _02989_ VGND VGND VPWR
+ VPWR _02990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09513_ _04528_ VGND VGND VPWR VPWR _00061_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06725_ u_rf.reg5_q\[6\] _01568_ _01555_ u_rf.reg6_q\[6\] _01982_ VGND VGND VPWR
+ VPWR _01983_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_121_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09444_ u_rf.reg2_q\[30\] _04490_ _04427_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__mux2_1
X_06656_ u_decod.pc_q_o\[2\] u_decod.pc_q_o\[3\] u_decod.pc_q_o\[4\] u_decod.pc_q_o\[5\]
+ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__and4_1
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09375_ u_decod.rf_ff_res_data_i\[8\] VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06587_ _01841_ _01850_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_613 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08326_ net475 _03259_ _03522_ _03340_ VGND VGND VPWR VPWR u_decod.rs1_data\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08257_ u_decod.exe_ff_res_data_i\[4\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[4\]
+ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__a221o_1
X_08188_ u_rf.reg6_q\[2\] _03387_ _03388_ u_rf.reg13_q\[2\] _03389_ VGND VGND VPWR
+ VPWR _03390_ sky130_fd_sc_hd__a221o_1
X_07208_ net40 net100 VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07139_ u_rf.reg29_q\[14\] _01628_ _01653_ u_rf.reg22_q\[14\] VGND VGND VPWR VPWR
+ _02381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_565 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10150_ _04886_ VGND VGND VPWR VPWR _00340_ sky130_fd_sc_hd__clkbuf_1
X_10081_ u_rf.reg9_q\[20\] _04469_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10983_ _05345_ VGND VGND VPWR VPWR _00714_ sky130_fd_sc_hd__clkbuf_1
X_12722_ clknet_leaf_40_clk _00759_ net279 VGND VGND VPWR VPWR u_rf.reg23_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ clknet_leaf_5_clk _00690_ net215 VGND VGND VPWR VPWR u_rf.reg21_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11604_ _04753_ u_rf.reg31_q\[15\] _05668_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__mux2_1
X_12584_ clknet_leaf_19_clk _00621_ net281 VGND VGND VPWR VPWR u_rf.reg19_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11535_ _05637_ VGND VGND VPWR VPWR _00974_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11466_ _04751_ u_rf.reg29_q\[14\] _05596_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11397_ _05564_ VGND VGND VPWR VPWR _00909_ sky130_fd_sc_hd__clkbuf_1
X_10417_ _05044_ VGND VGND VPWR VPWR _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _04724_ u_rf.reg13_q\[1\] _05006_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__mux2_1
X_10279_ _04961_ VGND VGND VPWR VPWR _00394_ sky130_fd_sc_hd__clkbuf_1
X_12018_ clknet_leaf_81_clk u_exe.bu_pc_res\[31\] net367 VGND VGND VPWR VPWR u_exe.pc_data_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_clk clknet_4_0_0_clk VGND VGND VPWR VPWR clknet_leaf_139_clk sky130_fd_sc_hd__clkbuf_16
X_06510_ _01674_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__buf_6
X_07490_ _01528_ _02695_ _02717_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06441_ net44 _01487_ _01488_ net41 _01709_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09160_ _04284_ _04286_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__nand2_1
X_06372_ _01641_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__buf_6
XFILLER_0_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09091_ _04226_ _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08111_ _03230_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_545 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08042_ u_decod.dec0.instr_i\[19\] _03172_ _03173_ VGND VGND VPWR VPWR _03248_ sky130_fd_sc_hd__and3_2
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_598 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09993_ u_rf.reg8_q\[11\] _04451_ _04801_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__mux2_1
X_08944_ _04042_ _04100_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__nor2_1
XFILLER_0_110_795 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ _03998_ _04041_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__nor2_1
X_07826_ u_decod.rf_ff_res_data_i\[28\] _02358_ _02743_ _03020_ _03039_ VGND VGND
+ VPWR VPWR _03040_ sky130_fd_sc_hd__a221o_1
X_07757_ u_decod.dec0.funct7\[2\] _01224_ _02646_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__a21o_1
X_06708_ _01506_ _01958_ _01966_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__a21oi_1
X_07688_ _02906_ _02907_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[25\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_32_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09427_ _04479_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06639_ _01895_ _01900_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[4\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_851 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09358_ u_rf.reg2_q\[2\] _04432_ _04428_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08309_ u_rf.reg9_q\[7\] _03348_ _03349_ u_rf.reg20_q\[7\] VGND VGND VPWR VPWR _03506_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11320_ _05523_ VGND VGND VPWR VPWR _00873_ sky130_fd_sc_hd__clkbuf_1
X_09289_ _04391_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_1
XFILLER_0_35_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11251_ u_rf.reg26_q\[9\] net471 _05477_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__mux2_1
X_10202_ _04914_ VGND VGND VPWR VPWR _00364_ sky130_fd_sc_hd__clkbuf_1
X_11182_ _05450_ VGND VGND VPWR VPWR _00808_ sky130_fd_sc_hd__clkbuf_1
X_10133_ _04877_ VGND VGND VPWR VPWR _00332_ sky130_fd_sc_hd__clkbuf_1
X_10064_ u_rf.reg9_q\[12\] _04453_ _04838_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_535 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10966_ _05336_ VGND VGND VPWR VPWR _00706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10897_ u_rf.reg21_q\[2\] _04943_ _05297_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__mux2_1
X_12705_ clknet_leaf_118_clk _00742_ net326 VGND VGND VPWR VPWR u_rf.reg23_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12636_ clknet_leaf_127_clk _00673_ net237 VGND VGND VPWR VPWR u_rf.reg21_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12567_ clknet_leaf_70_clk _00604_ net352 VGND VGND VPWR VPWR u_rf.reg18_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12498_ clknet_leaf_38_clk _00535_ net274 VGND VGND VPWR VPWR u_rf.reg16_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11518_ _05628_ VGND VGND VPWR VPWR _00966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11449_ _04734_ u_rf.reg29_q\[6\] _05585_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__mux2_1
X_06990_ u_decod.rs1_data_q\[27\] _01454_ _01753_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__o21a_1
X_05941_ _01223_ VGND VGND VPWR VPWR u_decod.dec0.is_shift sky130_fd_sc_hd__clkbuf_1
X_08660_ u_rf.reg31_q\[23\] _03504_ _03505_ u_rf.reg11_q\[23\] _03840_ VGND VGND VPWR
+ VPWR _03841_ sky130_fd_sc_hd__a221o_1
X_05872_ u_decod.pc0_q_i\[23\] _01168_ VGND VGND VPWR VPWR _01171_ sky130_fd_sc_hd__and2_4
XFILLER_0_89_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07611_ _02629_ _02833_ _01905_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__mux2_1
X_08591_ u_rf.reg18_q\[20\] _03262_ _03263_ u_rf.reg23_q\[20\] _03774_ VGND VGND VPWR
+ VPWR _03775_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_85_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07542_ _02765_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07473_ u_rf.reg9_q\[21\] _01636_ _01671_ u_rf.reg27_q\[21\] _02700_ VGND VGND VPWR
+ VPWR _02701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09212_ _04318_ _04320_ _04324_ _04323_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06424_ _01479_ _01689_ _01692_ _01441_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09143_ _04270_ _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06355_ _01624_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09074_ _04004_ _04207_ _04208_ _04213_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[2\]
+ sky130_fd_sc_hd__a2bb2o_1
X_06286_ _01555_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08025_ _03170_ _03173_ _03204_ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__and3_4
XFILLER_0_13_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09976_ u_rf.reg8_q\[3\] _04434_ _04790_ VGND VGND VPWR VPWR _04794_ sky130_fd_sc_hd__mux2_1
X_08927_ _04084_ _04085_ VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__nor2_2
X_08858_ u_decod.rs1_data_q\[4\] u_decod.branch_imm_q_o\[4\] _04026_ _04019_ VGND
+ VGND VPWR VPWR _04027_ sky130_fd_sc_hd__a31o_1
X_07809_ u_rf.reg25_q\[28\] _01783_ _02379_ u_rf.reg17_q\[28\] VGND VGND VPWR VPWR
+ _03023_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _03957_ _03959_ _03961_ _03963_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__or4_1
X_10820_ u_rf.reg19_q\[31\] _05003_ _05223_ VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10751_ _05221_ VGND VGND VPWR VPWR _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10682_ u_rf.reg17_q\[30\] _05001_ _05151_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12421_ clknet_leaf_122_clk _00458_ net241 VGND VGND VPWR VPWR u_rf.reg14_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12352_ clknet_leaf_114_clk _00389_ net323 VGND VGND VPWR VPWR u_rf.reg12_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12283_ clknet_leaf_13_clk _00320_ net243 VGND VGND VPWR VPWR u_rf.reg10_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11303_ _04724_ u_rf.reg27_q\[1\] _05513_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11234_ _05478_ VGND VGND VPWR VPWR _00832_ sky130_fd_sc_hd__clkbuf_1
X_11165_ u_rf.reg25_q\[0\] _04935_ _05441_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__mux2_1
X_11096_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__buf_6
X_10116_ _04868_ VGND VGND VPWR VPWR _00324_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10047_ u_rf.reg9_q\[4\] _04436_ _04827_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__mux2_1
Xhold80 u_decod.pc0_q_i\[19\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold91 u_decod.pc0_q_i\[9\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11998_ clknet_leaf_84_clk u_exe.bu_pc_res\[11\] net364 VGND VGND VPWR VPWR u_exe.pc_data_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10949_ u_rf.reg21_q\[27\] _04995_ _05319_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_760 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_849 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12619_ clknet_leaf_135_clk _00656_ net208 VGND VGND VPWR VPWR u_rf.reg20_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06140_ _01276_ _01278_ _01410_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_470 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06071_ _01301_ _01300_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_479 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _04700_ VGND VGND VPWR VPWR _00206_ sky130_fd_sc_hd__clkbuf_1
X_09761_ _04663_ VGND VGND VPWR VPWR _00174_ sky130_fd_sc_hd__clkbuf_1
X_06973_ u_rf.reg6_q\[11\] _01556_ _01622_ u_rf.reg24_q\[11\] _02220_ VGND VGND VPWR
+ VPWR _02221_ sky130_fd_sc_hd__a221o_1
X_08712_ u_rf.reg27_q\[25\] _03365_ _03320_ u_rf.reg19_q\[25\] VGND VGND VPWR VPWR
+ _03891_ sky130_fd_sc_hd__a22o_1
X_05924_ _01213_ VGND VGND VPWR VPWR u_decod.dec0.rd_v sky130_fd_sc_hd__clkbuf_2
X_09692_ _04625_ VGND VGND VPWR VPWR _00143_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer12 u_decod.pc0_q_i\[4\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_2
X_05855_ _01099_ _01156_ _01157_ _01158_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__a31o_1
X_08643_ u_rf.reg25_q\[22\] _03315_ _03328_ u_rf.reg12_q\[22\] _03824_ VGND VGND VPWR
+ VPWR _03825_ sky130_fd_sc_hd__a221o_1
Xrebuffer23 net398 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
Xrebuffer34 _04040_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05786_ _01098_ VGND VGND VPWR VPWR _01106_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08574_ u_rf.reg9_q\[19\] _03293_ _03295_ u_rf.reg20_q\[19\] VGND VGND VPWR VPWR
+ _03759_ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07525_ u_rf.reg7_q\[22\] _01562_ _02665_ u_rf.reg19_q\[22\] VGND VGND VPWR VPWR
+ _02751_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_321 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_61_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07456_ _01905_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07387_ _02446_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__buf_2
X_06407_ _01633_ _01647_ _01661_ _01676_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09126_ _04256_ _04257_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__and2_1
X_06338_ _01607_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_802 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09057_ u_decod.branch_imm_q_o\[0\] u_decod.pc_q_o\[0\] VGND VGND VPWR VPWR _04199_
+ sky130_fd_sc_hd__or2_1
X_06269_ u_decod.rf_ff_rd_adr_q_i\[4\] VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_446 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08008_ u_rf.reg9_q\[31\] _03212_ _03213_ u_rf.reg20_q\[31\] VGND VGND VPWR VPWR
+ _03214_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09959_ _04782_ u_rf.reg7_q\[29\] _04764_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12970_ clknet_leaf_27_clk _01007_ net259 VGND VGND VPWR VPWR u_rf.reg31_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_11921_ clknet_leaf_102_clk u_decod.rs1_data\[9\] net337 VGND VGND VPWR VPWR u_decod.rs1_data_q\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_142_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ clknet_leaf_29_clk _00079_ net257 VGND VGND VPWR VPWR u_rf.reg0_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10803_ _05249_ VGND VGND VPWR VPWR _00630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_clk clknet_4_13_0_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
X_11783_ clknet_leaf_84_clk net135 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_67_376 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10734_ u_rf.reg18_q\[22\] _04985_ _05210_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10665_ _05176_ VGND VGND VPWR VPWR _00565_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12404_ clknet_leaf_31_clk _00441_ net261 VGND VGND VPWR VPWR u_rf.reg13_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_711 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12335_ clknet_leaf_43_clk _00372_ net294 VGND VGND VPWR VPWR u_rf.reg11_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ u_rf.reg16_q\[21\] _04983_ _05138_ VGND VGND VPWR VPWR _05140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_654 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12266_ clknet_leaf_29_clk _00303_ net257 VGND VGND VPWR VPWR u_rf.reg9_q\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11217_ u_rf.reg25_q\[25\] _04991_ _05463_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__mux2_1
X_12197_ clknet_leaf_121_clk _00234_ net248 VGND VGND VPWR VPWR u_rf.reg7_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11148_ _05432_ VGND VGND VPWR VPWR _00792_ sky130_fd_sc_hd__clkbuf_1
X_11079_ _04772_ u_rf.reg23_q\[24\] _05391_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_33 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07310_ _02189_ _02499_ _02544_ _01505_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08290_ u_rf.reg26_q\[6\] _03203_ _03206_ u_rf.reg21_q\[6\] VGND VGND VPWR VPWR _03488_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07241_ u_rf.reg30_q\[16\] _01579_ _01591_ u_rf.reg18_q\[16\] VGND VGND VPWR VPWR
+ _02479_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07172_ _01291_ _02412_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06123_ _01288_ _01357_ _01393_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__nand3_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06054_ u_decod.rs2_data_q\[7\] u_decod.rs1_data_q\[7\] VGND VGND VPWR VPWR _01325_
+ sky130_fd_sc_hd__nor2_1
Xfanout304 net305 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_838 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout348 net373 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_2
Xfanout326 net327 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_4
X_09813_ _04691_ VGND VGND VPWR VPWR _00198_ sky130_fd_sc_hd__clkbuf_1
Xfanout315 net318 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__buf_2
Xfanout337 net338 VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__buf_2
Xfanout359 net373 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_2
X_09744_ _04654_ VGND VGND VPWR VPWR _00166_ sky130_fd_sc_hd__clkbuf_1
X_06956_ u_decod.dec0.instr_i\[20\] _01205_ _01241_ u_decod.dec0.instr_i\[7\] _02203_
+ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__a221o_2
X_06887_ _01949_ _01754_ _01950_ _02137_ _01450_ _01467_ VGND VGND VPWR VPWR _02138_
+ sky130_fd_sc_hd__mux4_1
X_09675_ _04616_ VGND VGND VPWR VPWR _00135_ sky130_fd_sc_hd__clkbuf_1
X_05907_ u_decod.dec0.funct3\[1\] _01077_ VGND VGND VPWR VPWR _01197_ sky130_fd_sc_hd__or2_1
X_08626_ u_rf.reg0_q\[21\] _03420_ _03421_ u_rf.reg12_q\[21\] _03808_ VGND VGND VPWR
+ VPWR _03809_ sky130_fd_sc_hd__a221o_1
X_05838_ _01143_ _01144_ _01145_ VGND VGND VPWR VPWR _01146_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_6_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
X_08557_ u_rf.reg9_q\[18\] _03293_ _03295_ u_rf.reg20_q\[18\] VGND VGND VPWR VPWR
+ _03743_ sky130_fd_sc_hd__a22o_1
X_05769_ u_decod.dec0.instr_i\[4\] _01087_ VGND VGND VPWR VPWR _01092_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08488_ u_rf.reg26_q\[15\] _03284_ _03345_ u_rf.reg21_q\[15\] VGND VGND VPWR VPWR
+ _03677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07508_ _02686_ _02734_ _01480_ VGND VGND VPWR VPWR _02735_ sky130_fd_sc_hd__mux2_1
X_07439_ _02657_ _02668_ _01680_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__o21a_2
XFILLER_0_64_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10450_ _05061_ VGND VGND VPWR VPWR _00465_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09109_ _04034_ _04207_ _04208_ _04243_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[7\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10381_ _04757_ u_rf.reg13_q\[17\] _05017_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_265 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12120_ clknet_leaf_65_clk _00157_ net346 VGND VGND VPWR VPWR u_rf.reg4_q\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12051_ clknet_leaf_91_clk u_decod.exe_ff_res_data_i\[31\] net344 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[31\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_2_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11002_ _05332_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_102_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_144_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ clknet_leaf_62_clk _00990_ net341 VGND VGND VPWR VPWR u_rf.reg30_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11904_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[25\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12884_ clknet_leaf_22_clk _00921_ net285 VGND VGND VPWR VPWR u_rf.reg28_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_337 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11835_ clknet_leaf_114_clk net24 net328 VGND VGND VPWR VPWR u_decod.dec0.funct7\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11766_ clknet_leaf_47_clk _00058_ net300 VGND VGND VPWR VPWR u_rf.reg1_q\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_562 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10717_ u_rf.reg18_q\[14\] _04968_ _05199_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11697_ _05723_ VGND VGND VPWR VPWR _01050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10648_ _05167_ VGND VGND VPWR VPWR _00557_ sky130_fd_sc_hd__clkbuf_1
Xrebuffer3 net376 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10579_ u_rf.reg16_q\[13\] _04966_ _05127_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12318_ clknet_leaf_123_clk _00355_ net241 VGND VGND VPWR VPWR u_rf.reg11_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_484 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12249_ clknet_leaf_62_clk _00286_ net343 VGND VGND VPWR VPWR u_rf.reg8_q\[30\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07790_ _01266_ _03003_ _02332_ VGND VGND VPWR VPWR _03005_ sky130_fd_sc_hd__o21a_1
X_06810_ u_rf.reg30_q\[8\] _01578_ _01623_ u_rf.reg28_q\[8\] VGND VGND VPWR VPWR _02064_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06741_ _01442_ _01997_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__nand2_1
X_09460_ u_rf.reg1_q\[4\] _04436_ _04496_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06672_ _01925_ _01927_ _01929_ _01931_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__or4_1
X_08411_ _03597_ _03599_ _03601_ _03603_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_35_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09391_ u_decod.rf_ff_res_data_i\[13\] VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_16_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08342_ u_rf.reg1_q\[8\] _03311_ _03313_ u_rf.reg14_q\[8\] VGND VGND VPWR VPWR _03538_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_157_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08273_ u_rf.reg24_q\[5\] _03302_ _03272_ u_rf.reg29_q\[5\] _03471_ VGND VGND VPWR
+ VPWR _03472_ sky130_fd_sc_hd__a221o_1
X_07224_ _01764_ _02461_ _02462_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__or3_2
XFILLER_0_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07155_ _02394_ _02396_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[14\] sky130_fd_sc_hd__xor2_1
XFILLER_0_15_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06106_ u_decod.rs2_data_q\[19\] _01376_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__or2_1
X_07086_ _02328_ _02329_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[13\] sky130_fd_sc_hd__xor2_1
XFILLER_0_30_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06037_ _01306_ _01307_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07988_ u_decod.rf_ff_rd_adr_q_i\[0\] u_decod.dec0.instr_i\[15\] VGND VGND VPWR VPWR
+ _03194_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09727_ _01534_ _04424_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__nor2_1
X_06939_ _01424_ _02139_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09658_ _04423_ _04606_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_2_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08609_ u_decod.exe_ff_res_data_i\[20\] _03669_ _03670_ u_decod.rf_ff_res_data_i\[20\]
+ _03792_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a221o_1
X_09589_ _04423_ _04569_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__nor2_4
X_11620_ _05682_ VGND VGND VPWR VPWR _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11551_ _04768_ u_rf.reg30_q\[22\] _05643_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_357 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10502_ _05077_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__buf_6
XFILLER_0_53_828 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11482_ _05609_ VGND VGND VPWR VPWR _00949_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10433_ _05052_ VGND VGND VPWR VPWR _00457_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10364_ _04740_ u_rf.reg13_q\[9\] _05006_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12103_ clknet_leaf_4_clk _00140_ net212 VGND VGND VPWR VPWR u_rf.reg4_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10295_ u_decod.rf_ff_res_data_i\[16\] VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__buf_2
XFILLER_0_109_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12034_ clknet_leaf_91_clk u_decod.exe_ff_res_data_i\[14\] net344 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[14\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_70_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_69_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12936_ clknet_leaf_58_clk _00973_ net291 VGND VGND VPWR VPWR u_rf.reg30_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_12867_ clknet_leaf_112_clk _00904_ net321 VGND VGND VPWR VPWR u_rf.reg28_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_157_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ clknet_leaf_105_clk net5 net319 VGND VGND VPWR VPWR u_decod.dec0.funct3\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12798_ clknet_leaf_123_clk _00835_ net241 VGND VGND VPWR VPWR u_rf.reg26_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11749_ clknet_leaf_108_clk _00041_ net312 VGND VGND VPWR VPWR u_rf.reg1_q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_119_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08960_ _04113_ VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__inv_2
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07911_ u_rf.reg24_q\[30\] _01784_ _02379_ u_rf.reg17_q\[30\] VGND VGND VPWR VPWR
+ _03121_ sky130_fd_sc_hd__a22o_1
X_08891_ u_decod.rs1_data_q\[11\] u_decod.branch_imm_q_o\[11\] VGND VGND VPWR VPWR
+ _04055_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_87_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07842_ _01443_ _03049_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_108_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07773_ u_rf.reg26_q\[27\] _02368_ _02385_ u_rf.reg20_q\[27\] VGND VGND VPWR VPWR
+ _02989_ sky130_fd_sc_hd__a22o_1
X_09512_ u_rf.reg1_q\[29\] _04488_ _04518_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06724_ u_rf.reg31_q\[6\] _01615_ _01648_ u_rf.reg4_q\[6\] VGND VGND VPWR VPWR _01982_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09443_ u_decod.rf_ff_res_data_i\[30\] VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__buf_2
X_06655_ _01058_ _01915_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09374_ _04443_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_96_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08325_ u_decod.exe_ff_res_data_i\[7\] _03260_ _03261_ u_decod.rf_ff_res_data_i\[7\]
+ _03521_ VGND VGND VPWR VPWR _03522_ sky130_fd_sc_hd__a221o_1
X_06586_ _01843_ _01845_ _01847_ _01849_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08256_ _03443_ _03455_ _03337_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08187_ u_rf.reg15_q\[2\] _03237_ _03238_ u_rf.reg24_q\[2\] VGND VGND VPWR VPWR _03389_
+ sky130_fd_sc_hd__a22o_1
X_07207_ u_decod.unsign_ext_q_o _02445_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_43_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07138_ _01791_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_883 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07069_ u_rf.reg31_q\[13\] _01615_ _01658_ u_rf.reg14_q\[13\] _02312_ VGND VGND VPWR
+ VPWR _02313_ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10080_ _04826_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_7_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10982_ u_rf.reg22_q\[10\] _04959_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__mux2_1
X_12721_ clknet_leaf_56_clk _00758_ net293 VGND VGND VPWR VPWR u_rf.reg23_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12652_ clknet_leaf_26_clk _00689_ net265 VGND VGND VPWR VPWR u_rf.reg21_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _05673_ VGND VGND VPWR VPWR _01006_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_474 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12583_ clknet_leaf_4_clk _00620_ net214 VGND VGND VPWR VPWR u_rf.reg19_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11534_ _04751_ u_rf.reg30_q\[14\] _05632_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_152_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11465_ _05600_ VGND VGND VPWR VPWR _00941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10416_ _04724_ u_rf.reg14_q\[1\] _05042_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__mux2_1
X_11396_ u_rf.reg28_q\[13\] u_decod.rf_ff_res_data_i\[13\] _05560_ VGND VGND VPWR
+ VPWR _05564_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_405 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10347_ _05007_ VGND VGND VPWR VPWR _00416_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ u_rf.reg12_q\[10\] _04959_ _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12017_ clknet_leaf_81_clk u_exe.bu_pc_res\[30\] net368 VGND VGND VPWR VPWR u_exe.pc_data_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_12919_ clknet_leaf_71_clk _00956_ net354 VGND VGND VPWR VPWR u_rf.reg29_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06440_ net64 _01489_ _01490_ net50 VGND VGND VPWR VPWR _01709_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_516 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06371_ _01640_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_145_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09090_ u_decod.pc_q_o\[5\] u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _04227_
+ sky130_fd_sc_hd__and2_1
X_08110_ _03229_ VGND VGND VPWR VPWR _03314_ sky130_fd_sc_hd__buf_6
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08041_ _03188_ _03173_ _03209_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__and3_4
XFILLER_0_43_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_557 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_741 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09992_ _04802_ VGND VGND VPWR VPWR _00266_ sky130_fd_sc_hd__clkbuf_1
X_08943_ _04096_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_4_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08874_ _04037_ net408 VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__xnor2_1
X_07825_ _03029_ _03038_ _02359_ VGND VGND VPWR VPWR _03039_ sky130_fd_sc_hd__o21a_1
X_07756_ _02972_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[27\] sky130_fd_sc_hd__inv_2
X_06707_ _01058_ _01960_ _01965_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__a21o_1
X_09426_ u_rf.reg2_q\[24\] _04478_ _04470_ VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__mux2_1
X_07687_ _02862_ _02864_ net200 VGND VGND VPWR VPWR _02907_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06638_ _01897_ _01899_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__nand2_1
X_09357_ u_decod.rf_ff_res_data_i\[2\] VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06569_ u_rf.reg25_q\[3\] _01575_ _01641_ u_rf.reg26_q\[3\] VGND VGND VPWR VPWR _01833_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08308_ _03291_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__buf_8
XFILLER_0_90_731 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _04385_ u_decod.rs2_data_q\[7\] _04386_ VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__and3_1
XFILLER_0_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08239_ u_rf.reg26_q\[4\] _03284_ _03286_ u_rf.reg21_q\[4\] VGND VGND VPWR VPWR _03439_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11250_ _05486_ VGND VGND VPWR VPWR _00840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10201_ _04747_ u_rf.reg11_q\[12\] _04911_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__mux2_1
X_11181_ u_rf.reg25_q\[8\] _04955_ _05441_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10132_ u_rf.reg10_q\[12\] _04453_ _04874_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__mux2_1
X_10063_ _04840_ VGND VGND VPWR VPWR _00299_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10965_ u_rf.reg22_q\[2\] _04943_ _05333_ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__mux2_1
X_12704_ clknet_leaf_117_clk _00741_ net327 VGND VGND VPWR VPWR u_rf.reg23_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10896_ _05299_ VGND VGND VPWR VPWR _00673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12635_ clknet_leaf_122_clk _00672_ net242 VGND VGND VPWR VPWR u_rf.reg21_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12566_ clknet_leaf_49_clk _00603_ net308 VGND VGND VPWR VPWR u_rf.reg18_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11517_ _04734_ u_rf.reg30_q\[6\] _05621_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12497_ clknet_leaf_53_clk _00534_ net302 VGND VGND VPWR VPWR u_rf.reg16_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11448_ _05591_ VGND VGND VPWR VPWR _00933_ sky130_fd_sc_hd__clkbuf_1
X_11379_ u_rf.reg28_q\[5\] u_decod.rf_ff_res_data_i\[5\] _05549_ VGND VGND VPWR VPWR
+ _05555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05940_ _01220_ _01222_ VGND VGND VPWR VPWR _01223_ sky130_fd_sc_hd__or2_1
X_05871_ net481 _01142_ _01132_ net79 _01170_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__a221o_1
XFILLER_0_56_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08590_ u_rf.reg4_q\[20\] _03264_ _03266_ u_rf.reg17_q\[20\] VGND VGND VPWR VPWR
+ _03774_ sky130_fd_sc_hd__a22o_1
X_07610_ u_decod.rs1_data_q\[24\] _01388_ u_decod.rs1_data_q\[8\] _01061_ _01467_
+ _01461_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__mux4_1
X_07541_ _02089_ _02487_ _02672_ _02766_ net200 VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__a41o_1
XFILLER_0_89_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07472_ u_rf.reg12_q\[21\] _01609_ _01673_ u_rf.reg2_q\[21\] VGND VGND VPWR VPWR
+ _02700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09211_ _04318_ _04320_ _04324_ _04330_ _04323_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__a311o_1
XFILLER_0_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06423_ _01690_ _01691_ _01422_ VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09142_ _04265_ _04260_ _04262_ _04263_ _04271_ VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06354_ _01623_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__buf_6
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_866 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09073_ _04209_ _04212_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06285_ _01554_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__buf_6
XFILLER_0_130_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08024_ _03188_ _03201_ _03204_ VGND VGND VPWR VPWR _03230_ sky130_fd_sc_hd__and3_2
XFILLER_0_13_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09975_ _04793_ VGND VGND VPWR VPWR _00258_ sky130_fd_sc_hd__clkbuf_1
X_08926_ _01388_ u_decod.branch_imm_q_o\[16\] VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__and2_1
XFILLER_0_99_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08857_ u_decod.rs1_data_q\[5\] u_decod.branch_imm_q_o\[5\] VGND VGND VPWR VPWR _04026_
+ sky130_fd_sc_hd__or2_1
X_07808_ u_rf.reg21_q\[28\] _02364_ _01776_ u_rf.reg2_q\[28\] _03021_ VGND VGND VPWR
+ VPWR _03022_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_28_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ u_rf.reg25_q\[29\] _03370_ _03313_ u_rf.reg14_q\[29\] _03962_ VGND VGND VPWR
+ VPWR _03963_ sky130_fd_sc_hd__a221o_1
X_07739_ _01283_ _01409_ _02911_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__or3b_1
XFILLER_0_95_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10750_ u_rf.reg18_q\[30\] _05001_ _05187_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_867 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10681_ _05184_ VGND VGND VPWR VPWR _00573_ sky130_fd_sc_hd__clkbuf_1
X_09409_ u_decod.rf_ff_res_data_i\[19\] VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__buf_2
XFILLER_0_36_901 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_260 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12420_ clknet_leaf_109_clk _00457_ net313 VGND VGND VPWR VPWR u_rf.reg14_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_466 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12351_ clknet_leaf_132_clk _00388_ net228 VGND VGND VPWR VPWR u_rf.reg12_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12282_ clknet_leaf_61_clk _00319_ net339 VGND VGND VPWR VPWR u_rf.reg9_q\[31\] sky130_fd_sc_hd__dfrtp_1
X_11302_ _05514_ VGND VGND VPWR VPWR _00864_ sky130_fd_sc_hd__clkbuf_1
X_11233_ u_rf.reg26_q\[0\] net503 _05477_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__mux2_1
X_11164_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_147_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11095_ _04788_ _05114_ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__nor2_4
X_10115_ u_rf.reg10_q\[4\] _04436_ _04863_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10046_ _04831_ VGND VGND VPWR VPWR _00291_ sky130_fd_sc_hd__clkbuf_1
Xhold81 u_decod.pc0_q_i\[25\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold70 u_decod.pc0_q_i\[14\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 u_decod.dec0.instr_i\[3\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_133_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11997_ clknet_leaf_84_clk u_exe.bu_pc_res\[10\] net364 VGND VGND VPWR VPWR u_exe.pc_data_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10948_ _05326_ VGND VGND VPWR VPWR _00698_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_772 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10879_ _05289_ VGND VGND VPWR VPWR _00666_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12618_ clknet_leaf_30_clk _00655_ net262 VGND VGND VPWR VPWR u_rf.reg20_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_293 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12549_ clknet_leaf_111_clk _00586_ net316 VGND VGND VPWR VPWR u_rf.reg18_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_1 _01099_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06070_ _01332_ _01336_ _01337_ _01340_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09760_ u_rf.reg5_q\[14\] _04457_ _04658_ VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__mux2_1
X_06972_ u_rf.reg15_q\[11\] _01600_ _01612_ u_rf.reg23_q\[11\] VGND VGND VPWR VPWR
+ _02220_ sky130_fd_sc_hd__a22o_1
X_08711_ u_rf.reg0_q\[25\] _03420_ _03421_ u_rf.reg12_q\[25\] _03889_ VGND VGND VPWR
+ VPWR _03890_ sky130_fd_sc_hd__a221o_1
X_09691_ u_rf.reg4_q\[15\] _04459_ _04619_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__mux2_1
X_05923_ _01204_ _01208_ _01212_ VGND VGND VPWR VPWR _01213_ sky130_fd_sc_hd__or3b_1
X_08642_ u_rf.reg0_q\[22\] _03174_ _03238_ u_rf.reg24_q\[22\] VGND VGND VPWR VPWR
+ _03824_ sky130_fd_sc_hd__a22o_1
X_05854_ net515 _01118_ _01119_ net74 VGND VGND VPWR VPWR _01158_ sky130_fd_sc_hd__a22o_1
Xrebuffer24 net399 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
Xrebuffer13 _04053_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer35 u_decod.rs1_data_q\[1\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_1
XFILLER_0_107_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05785_ _01104_ VGND VGND VPWR VPWR _01105_ sky130_fd_sc_hd__clkbuf_4
X_08573_ u_rf.reg8_q\[19\] _03270_ _03272_ u_rf.reg29_q\[19\] _03757_ VGND VGND VPWR
+ VPWR _03758_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_402 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07524_ u_rf.reg14_q\[22\] _02367_ _01654_ u_rf.reg22_q\[22\] _02749_ VGND VGND VPWR
+ VPWR _02750_ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_333 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07455_ _01358_ u_decod.rs1_data_q\[13\] u_decod.rs1_data_q\[5\] _01747_ _01468_
+ _01461_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06406_ u_rf.reg0_q\[0\] _01664_ _01668_ u_rf.reg8_q\[0\] _01675_ VGND VGND VPWR
+ VPWR _01676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07386_ _02616_ _02617_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[19\] sky130_fd_sc_hd__xor2_1
XFILLER_0_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09125_ u_decod.pc_q_o\[10\] u_decod.branch_imm_q_o\[10\] VGND VGND VPWR VPWR _04257_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06337_ _01513_ _01514_ _01577_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_131_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_814 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09056_ u_decod.branch_imm_q_o\[0\] u_decod.pc_q_o\[0\] VGND VGND VPWR VPWR _04198_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06268_ u_decod.dec0.instr_i\[24\] VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__buf_2
XFILLER_0_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08007_ u_decod.dec0.instr_i\[19\] _03172_ _03205_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__and3_4
X_06199_ _01061_ _01388_ u_decod.rs1_data_q\[8\] u_decod.rs1_data_q\[24\] _01466_
+ _01469_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__mux4_1
X_09958_ u_decod.rf_ff_res_data_i\[29\] VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _04069_ _04070_ VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09889_ _04735_ VGND VGND VPWR VPWR _00230_ sky130_fd_sc_hd__clkbuf_1
X_11920_ clknet_leaf_102_clk u_decod.rs1_data\[8\] net337 VGND VGND VPWR VPWR u_decod.rs1_data_q\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_142_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ clknet_leaf_20_clk _00078_ net280 VGND VGND VPWR VPWR u_rf.reg0_q\[14\] sky130_fd_sc_hd__dfrtp_1
X_10802_ u_rf.reg19_q\[22\] _04985_ _05246_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__mux2_1
X_11782_ clknet_leaf_85_clk net165 net364 VGND VGND VPWR VPWR u_decod.pc0_q_i\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10733_ _05212_ VGND VGND VPWR VPWR _00597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_826 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_709 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10664_ u_rf.reg17_q\[21\] _04983_ _05174_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10595_ _05139_ VGND VGND VPWR VPWR _00532_ sky130_fd_sc_hd__clkbuf_1
X_12403_ clknet_leaf_53_clk _00440_ net302 VGND VGND VPWR VPWR u_rf.reg13_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_408 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12334_ clknet_leaf_7_clk _00371_ net258 VGND VGND VPWR VPWR u_rf.reg11_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12265_ clknet_leaf_21_clk _00302_ net280 VGND VGND VPWR VPWR u_rf.reg9_q\[14\] sky130_fd_sc_hd__dfrtp_1
X_11216_ _05468_ VGND VGND VPWR VPWR _00824_ sky130_fd_sc_hd__clkbuf_1
X_12196_ clknet_leaf_109_clk _00233_ net313 VGND VGND VPWR VPWR u_rf.reg7_q\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11147_ u_rf.reg24_q\[24\] _04989_ _05427_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11078_ _05395_ VGND VGND VPWR VPWR _00759_ sky130_fd_sc_hd__clkbuf_1
X_10029_ _04821_ VGND VGND VPWR VPWR _00284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07240_ u_rf.reg20_q\[16\] _01644_ _01670_ u_rf.reg27_q\[16\] _02477_ VGND VGND VPWR
+ VPWR _02478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07171_ _02411_ _01435_ _01432_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_669 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06122_ _01375_ _01392_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06053_ _01322_ _01323_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__and2_1
Xfanout305 net310 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__buf_2
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09812_ u_rf.reg6_q\[6\] _04440_ _04684_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__mux2_1
Xfanout316 net318 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_4
Xfanout338 net374 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_4
Xfanout327 net334 VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__buf_4
Xfanout349 net359 VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09743_ u_rf.reg5_q\[6\] _04440_ _04647_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__mux2_1
X_06955_ _01227_ _01530_ u_decod.dec0.funct7\[6\] VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_05906_ net500 _01118_ _01119_ net89 _01196_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__a221o_1
XFILLER_0_69_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06886_ u_decod.rs1_data_q\[25\] _01454_ _02136_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__o21a_1
X_09674_ u_rf.reg4_q\[7\] _04442_ _04608_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__mux2_1
X_08625_ u_rf.reg28_q\[21\] _03556_ _03557_ u_rf.reg2_q\[21\] VGND VGND VPWR VPWR
+ _03808_ sky130_fd_sc_hd__a22o_1
X_05837_ u_decod.pc0_q_i\[14\] _01139_ VGND VGND VPWR VPWR _01145_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ u_rf.reg1_q\[18\] _03446_ _03332_ u_rf.reg2_q\[18\] _03741_ VGND VGND VPWR
+ VPWR _03742_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07507_ _02630_ _02733_ _01476_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__mux2_1
X_05768_ u_decod.dec0.instr_i\[0\] u_decod.dec0.funct3\[1\] u_decod.dec0.funct3\[2\]
+ VGND VGND VPWR VPWR _01091_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08487_ u_rf.reg31_q\[15\] _03504_ _03505_ u_rf.reg11_q\[15\] _03675_ VGND VGND VPWR
+ VPWR _03676_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07438_ _02659_ _02661_ _02663_ _02667_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07369_ u_rf.reg11_q\[19\] _01583_ _01642_ u_rf.reg26_q\[19\] VGND VGND VPWR VPWR
+ _02601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09108_ _04240_ _04242_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_482 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10380_ _05024_ VGND VGND VPWR VPWR _00432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09039_ _01280_ _01283_ _01361_ _01374_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__or4b_1
XFILLER_0_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12050_ clknet_leaf_90_clk u_decod.exe_ff_res_data_i\[30\] net346 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11001_ _05354_ VGND VGND VPWR VPWR _00723_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ clknet_leaf_67_clk _00989_ net349 VGND VGND VPWR VPWR u_rf.reg30_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_116_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11903_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[24\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_266 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12883_ clknet_leaf_66_clk _00920_ net356 VGND VGND VPWR VPWR u_rf.reg28_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_349 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11834_ clknet_leaf_104_clk net22 net322 VGND VGND VPWR VPWR u_decod.dec0.funct7\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_138_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11765_ clknet_leaf_32_clk _00057_ net263 VGND VGND VPWR VPWR u_rf.reg1_q\[25\] sky130_fd_sc_hd__dfrtp_1
X_11696_ u_decod.branch_imm_q_o\[26\] _02930_ _05717_ VGND VGND VPWR VPWR _05723_
+ sky130_fd_sc_hd__mux2_1
X_10716_ _05203_ VGND VGND VPWR VPWR _00589_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10647_ u_rf.reg17_q\[13\] _04966_ _05163_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 _04089_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_125_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10578_ _05130_ VGND VGND VPWR VPWR _00524_ sky130_fd_sc_hd__clkbuf_1
X_12317_ clknet_leaf_16_clk _00354_ net250 VGND VGND VPWR VPWR u_rf.reg11_q\[2\] sky130_fd_sc_hd__dfrtp_1
X_12248_ clknet_leaf_57_clk _00285_ net302 VGND VGND VPWR VPWR u_rf.reg8_q\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12179_ clknet_leaf_53_clk _00216_ net302 VGND VGND VPWR VPWR u_rf.reg6_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06740_ _01952_ _01996_ _01423_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__mux2_1
X_06671_ u_rf.reg18_q\[5\] _01591_ _01612_ u_rf.reg23_q\[5\] _01930_ VGND VGND VPWR
+ VPWR _01931_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_106_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08410_ u_rf.reg0_q\[11\] _03176_ _03329_ u_rf.reg12_q\[11\] _03602_ VGND VGND VPWR
+ VPWR _03603_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09390_ _04454_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_528 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08341_ u_rf.reg15_q\[8\] _03301_ _03303_ u_rf.reg24_q\[8\] _03536_ VGND VGND VPWR
+ VPWR _03537_ sky130_fd_sc_hd__a221o_1
X_08272_ u_rf.reg7_q\[5\] _03229_ _03230_ u_rf.reg25_q\[5\] VGND VGND VPWR VPWR _03471_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07223_ u_decod.pc_q_o\[15\] _02335_ u_decod.pc_q_o\[16\] VGND VGND VPWR VPWR _02462_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07154_ _02089_ _02395_ net201 VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06105_ u_decod.rs1_data_q\[19\] VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__buf_4
X_07085_ net199 _02278_ _02280_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06036_ u_decod.rs2_data_q\[8\] u_decod.rs1_data_q\[8\] VGND VGND VPWR VPWR _01307_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07987_ u_decod.rf_ff_rd_adr_q_i\[1\] _03190_ _03191_ _01536_ _03192_ VGND VGND VPWR
+ VPWR _03193_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ _01539_ u_decod.rf_write_v_q_i VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__and2_1
X_06938_ _01301_ _01820_ _02182_ _02186_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__o211ai_1
XTAP_TAPCELL_ROW_2_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09657_ u_decod.rf_ff_rd_adr_q_i\[0\] _04424_ _01532_ _01536_ VGND VGND VPWR VPWR
+ _04606_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_2_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06869_ u_rf.reg16_q\[9\] _01563_ _01629_ u_rf.reg17_q\[9\] VGND VGND VPWR VPWR _02121_
+ sky130_fd_sc_hd__a22o_1
X_08608_ _03782_ _03791_ _03378_ VGND VGND VPWR VPWR _03792_ sky130_fd_sc_hd__o21a_2
X_09588_ _01531_ _01536_ _04568_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__or3_4
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08539_ u_rf.reg16_q\[17\] _03248_ _03249_ u_rf.reg5_q\[17\] VGND VGND VPWR VPWR
+ _03726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_314 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11550_ _05645_ VGND VGND VPWR VPWR _00981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_453 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10501_ _05088_ VGND VGND VPWR VPWR _00489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_369 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11481_ _04766_ u_rf.reg29_q\[21\] _05607_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10432_ _04740_ u_rf.reg14_q\[9\] _05042_ VGND VGND VPWR VPWR _05052_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10363_ _05015_ VGND VGND VPWR VPWR _00424_ sky130_fd_sc_hd__clkbuf_1
X_12102_ clknet_leaf_139_clk _00139_ net202 VGND VGND VPWR VPWR u_rf.reg4_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ _04971_ VGND VGND VPWR VPWR _00399_ sky130_fd_sc_hd__clkbuf_1
X_12033_ clknet_leaf_93_clk u_decod.exe_ff_res_data_i\[13\] net344 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_57_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12935_ clknet_leaf_2_clk _00972_ net214 VGND VGND VPWR VPWR u_rf.reg30_q\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12866_ clknet_leaf_124_clk _00903_ net239 VGND VGND VPWR VPWR u_rf.reg28_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11817_ clknet_leaf_105_clk net4 net319 VGND VGND VPWR VPWR u_decod.dec0.funct3\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_141_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12797_ clknet_leaf_16_clk _00834_ net250 VGND VGND VPWR VPWR u_rf.reg26_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11748_ clknet_leaf_108_clk _00040_ net312 VGND VGND VPWR VPWR u_rf.reg1_q\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11679_ u_decod.branch_imm_q_o\[18\] _02551_ _05696_ VGND VGND VPWR VPWR _05714_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_290 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07910_ u_rf.reg9_q\[30\] _02360_ _01776_ u_rf.reg2_q\[30\] _03119_ VGND VGND VPWR
+ VPWR _03120_ sky130_fd_sc_hd__a221o_1
X_08890_ _04042_ _04054_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__nor2_1
XFILLER_0_20_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07841_ net133 _03050_ _03053_ _01746_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__a22o_1
X_07772_ u_rf.reg29_q\[27\] _01780_ _02364_ u_rf.reg21_q\[27\] _02987_ VGND VGND VPWR
+ VPWR _02988_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ _04527_ VGND VGND VPWR VPWR _00060_ sky130_fd_sc_hd__clkbuf_1
X_06723_ u_rf.reg0_q\[6\] _01662_ _01627_ u_rf.reg29_q\[6\] _01980_ VGND VGND VPWR
+ VPWR _01981_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09442_ _04489_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_121_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06654_ net60 _01487_ _01488_ net46 _01914_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09373_ u_rf.reg2_q\[7\] _04442_ _04428_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__mux2_1
X_06585_ u_rf.reg1_q\[3\] _01587_ _01625_ u_rf.reg28_q\[3\] _01848_ VGND VGND VPWR
+ VPWR _01849_ sky130_fd_sc_hd__a221o_1
XFILLER_0_148_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_319 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08324_ _03510_ _03520_ _03337_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__o21a_1
XFILLER_0_145_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_659 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08255_ _03445_ _03449_ _03452_ _03454_ VGND VGND VPWR VPWR _03455_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08186_ _03306_ VGND VGND VPWR VPWR _03388_ sky130_fd_sc_hd__buf_8
X_07206_ net98 net62 net57 _02049_ _02444_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_797 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07137_ _01631_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__buf_6
XFILLER_0_132_547 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07068_ u_rf.reg7_q\[13\] _01560_ _01641_ u_rf.reg26_q\[13\] VGND VGND VPWR VPWR
+ _02312_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06019_ u_decod.rs2_data_q\[15\] _01289_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_7_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09709_ _04634_ VGND VGND VPWR VPWR _00151_ sky130_fd_sc_hd__clkbuf_1
X_10981_ _05332_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__buf_6
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12720_ clknet_leaf_34_clk _00757_ net268 VGND VGND VPWR VPWR u_rf.reg23_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ clknet_leaf_1_clk _00688_ net223 VGND VGND VPWR VPWR u_rf.reg21_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _04751_ u_rf.reg31_q\[14\] _05668_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_842 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12582_ clknet_leaf_140_clk _00619_ net204 VGND VGND VPWR VPWR u_rf.reg19_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11533_ _05636_ VGND VGND VPWR VPWR _00973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_486 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_152_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _04749_ u_rf.reg29_q\[13\] _05596_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10415_ _05043_ VGND VGND VPWR VPWR _00448_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11395_ _05563_ VGND VGND VPWR VPWR _00908_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _04719_ u_rf.reg13_q\[0\] _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_567 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10277_ _04938_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_72_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12016_ clknet_leaf_81_clk u_exe.bu_pc_res\[29\] net368 VGND VGND VPWR VPWR u_exe.pc_data_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12918_ clknet_leaf_49_clk _00955_ net309 VGND VGND VPWR VPWR u_rf.reg29_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12849_ clknet_leaf_55_clk _00886_ net294 VGND VGND VPWR VPWR u_rf.reg27_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_144 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06370_ _01538_ _01553_ _01573_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08040_ _03188_ _03201_ _03209_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__and3_4
XFILLER_0_9_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_569 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09991_ u_rf.reg8_q\[10\] _04448_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__mux2_1
X_08942_ _04086_ _04089_ _04091_ _04098_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_110_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ _04025_ _04028_ _04032_ _04039_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07824_ _03031_ _03033_ _03035_ _03037_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07755_ _02332_ _02955_ _02956_ _02971_ VGND VGND VPWR VPWR _02972_ sky130_fd_sc_hd__a31oi_2
X_07686_ _02357_ u_decod.exe_ff_res_data_i\[25\] _02905_ VGND VGND VPWR VPWR _02906_
+ sky130_fd_sc_hd__a21oi_1
X_06706_ _01961_ _01431_ _01434_ _01330_ _01964_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__a221o_1
X_09425_ u_decod.rf_ff_res_data_i\[24\] VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_504 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06637_ _01804_ _01898_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06568_ u_decod.rf_ff_res_data_i\[3\] _01549_ _01773_ _01831_ VGND VGND VPWR VPWR
+ _01832_ sky130_fd_sc_hd__a22o_1
X_09356_ _04431_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08307_ _03289_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__buf_8
XFILLER_0_117_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06499_ _01313_ _01317_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09287_ _04390_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_1
XFILLER_0_90_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08238_ u_rf.reg8_q\[4\] _03271_ _03273_ u_rf.reg29_q\[4\] _03437_ VGND VGND VPWR
+ VPWR _03438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_134_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10200_ _04913_ VGND VGND VPWR VPWR _00363_ sky130_fd_sc_hd__clkbuf_1
X_08169_ u_rf.reg7_q\[1\] _03369_ _03370_ u_rf.reg25_q\[1\] _03371_ VGND VGND VPWR
+ VPWR _03372_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11180_ _05449_ VGND VGND VPWR VPWR _00807_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10131_ _04876_ VGND VGND VPWR VPWR _00331_ sky130_fd_sc_hd__clkbuf_1
X_10062_ u_rf.reg9_q\[11\] _04451_ _04838_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12703_ clknet_leaf_131_clk _00740_ net228 VGND VGND VPWR VPWR u_rf.reg23_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ _05335_ VGND VGND VPWR VPWR _00705_ sky130_fd_sc_hd__clkbuf_1
X_10895_ u_rf.reg21_q\[1\] _04941_ _05297_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__mux2_1
X_12634_ clknet_leaf_61_clk _00671_ net339 VGND VGND VPWR VPWR u_rf.reg20_q\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12565_ clknet_leaf_46_clk _00602_ net299 VGND VGND VPWR VPWR u_rf.reg18_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_341 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11516_ _05627_ VGND VGND VPWR VPWR _00965_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_653 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12496_ clknet_leaf_32_clk _00533_ net263 VGND VGND VPWR VPWR u_rf.reg16_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_697 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_889 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11447_ _04732_ u_rf.reg29_q\[5\] _05585_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_225 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11378_ _05554_ VGND VGND VPWR VPWR _00900_ sky130_fd_sc_hd__clkbuf_1
X_10329_ u_decod.rf_ff_res_data_i\[27\] VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__buf_2
XFILLER_0_147_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05870_ _01168_ _01144_ _01169_ VGND VGND VPWR VPWR _01170_ sky130_fd_sc_hd__and3b_1
XFILLER_0_89_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07540_ _02671_ _02718_ VGND VGND VPWR VPWR _02766_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07471_ u_rf.reg31_q\[21\] _01777_ _02697_ u_rf.reg4_q\[21\] _02698_ VGND VGND VPWR
+ VPWR _02699_ sky130_fd_sc_hd__a221o_1
X_09210_ _04328_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06422_ _01493_ _01459_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_604 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09141_ _04262_ u_decod.branch_imm_q_o\[10\] u_decod.pc_q_o\[10\] VGND VGND VPWR
+ VPWR _04271_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06353_ _01538_ _01514_ _01577_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__and3_2
XFILLER_0_115_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09072_ _04210_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08023_ _03171_ _03209_ _03205_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__and3_2
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06284_ _01512_ _01551_ _01553_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__and3_4
XTAP_TAPCELL_ROW_116_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_878 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09974_ u_rf.reg8_q\[2\] _04432_ _04790_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08925_ _01388_ u_decod.branch_imm_q_o\[16\] VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08856_ _04023_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__nor2_1
X_07807_ u_rf.reg10_q\[28\] _02380_ _02386_ u_rf.reg27_q\[28\] VGND VGND VPWR VPWR
+ _03021_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08787_ u_rf.reg24_q\[29\] _03302_ _03314_ u_rf.reg7_q\[29\] VGND VGND VPWR VPWR
+ _03962_ sky130_fd_sc_hd__a22o_1
X_05999_ _01268_ _01269_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__nor2_1
X_07738_ _01285_ _02911_ _01283_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__a21bo_1
X_07669_ u_rf.reg26_q\[25\] _01641_ _01649_ u_rf.reg4_q\[25\] VGND VGND VPWR VPWR
+ _02889_ sky130_fd_sc_hd__a22o_1
X_10680_ u_rf.reg17_q\[29\] _04999_ _05174_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09408_ _04466_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09339_ _04418_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__buf_1
XFILLER_0_63_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_881 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12350_ clknet_leaf_123_clk _00387_ net231 VGND VGND VPWR VPWR u_rf.reg12_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12281_ clknet_leaf_63_clk _00318_ net341 VGND VGND VPWR VPWR u_rf.reg9_q\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11301_ _04719_ u_rf.reg27_q\[0\] _05513_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11232_ _05476_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__buf_6
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_347 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11163_ _04644_ _04825_ _05295_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__and3_4
XFILLER_0_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10114_ _04867_ VGND VGND VPWR VPWR _00323_ sky130_fd_sc_hd__clkbuf_1
X_11094_ _05403_ VGND VGND VPWR VPWR _00767_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10045_ u_rf.reg9_q\[3\] _04434_ _04827_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__mux2_1
Xhold82 u_decod.pc0_q_i\[28\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 u_decod.pc0_q_i\[20\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold93 u_exe.pc_data_q\[9\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11996_ clknet_leaf_85_clk u_exe.bu_pc_res\[9\] net363 VGND VGND VPWR VPWR u_exe.pc_data_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10947_ u_rf.reg21_q\[26\] _04993_ _05319_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_47 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10878_ u_rf.reg20_q\[26\] _04993_ _05282_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__mux2_1
X_12617_ clknet_leaf_22_clk _00654_ net284 VGND VGND VPWR VPWR u_rf.reg20_q\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_54_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_620 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12548_ clknet_leaf_105_clk _00585_ net321 VGND VGND VPWR VPWR u_rf.reg18_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12479_ clknet_leaf_137_clk _00516_ net205 VGND VGND VPWR VPWR u_rf.reg16_q\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_2 _01206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ u_rf.reg20_q\[11\] _01645_ _01674_ u_rf.reg2_q\[11\] _02218_ VGND VGND VPWR
+ VPWR _02219_ sky130_fd_sc_hd__a221o_1
X_08710_ u_rf.reg28_q\[25\] _03330_ _03557_ u_rf.reg2_q\[25\] VGND VGND VPWR VPWR
+ _03889_ sky130_fd_sc_hd__a22o_1
X_09690_ _04624_ VGND VGND VPWR VPWR _00142_ sky130_fd_sc_hd__clkbuf_1
X_05922_ u_decod.dec0.instr_i\[0\] _01080_ _01075_ _01211_ VGND VGND VPWR VPWR _01212_
+ sky130_fd_sc_hd__nand4_1
X_05853_ u_decod.pc0_q_i\[18\] _01153_ VGND VGND VPWR VPWR _01157_ sky130_fd_sc_hd__nand2_1
X_08641_ _03816_ _03818_ _03820_ _03822_ VGND VGND VPWR VPWR _03823_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer25 net400 VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_1
Xrebuffer36 _01124_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer14 _04053_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
X_05784_ u_decod.flush_v net361 VGND VGND VPWR VPWR _01104_ sky130_fd_sc_hd__and2_1
X_08572_ u_rf.reg22_q\[19\] _03274_ _03276_ u_rf.reg3_q\[19\] VGND VGND VPWR VPWR
+ _03757_ sky130_fd_sc_hd__a22o_1
X_07523_ u_rf.reg15_q\[22\] _01601_ _02385_ u_rf.reg20_q\[22\] VGND VGND VPWR VPWR
+ _02749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07454_ _02625_ _02682_ _01425_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06405_ u_rf.reg27_q\[0\] _01671_ _01674_ u_rf.reg2_q\[0\] VGND VGND VPWR VPWR _01675_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_570 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_277 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07385_ _02489_ _02572_ _02573_ net199 VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_743 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06336_ _01605_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__buf_6
XFILLER_0_115_631 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09124_ u_decod.pc_q_o\[10\] u_decod.branch_imm_q_o\[10\] VGND VGND VPWR VPWR _04256_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_60_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_253 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ _04196_ VGND VGND VPWR VPWR _04197_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06267_ u_decod.dec0.instr_i\[23\] VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08006_ _03170_ _03201_ _03204_ VGND VGND VPWR VPWR _03212_ sky130_fd_sc_hd__and3_4
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_678 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06198_ _01468_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_481 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09957_ _04781_ VGND VGND VPWR VPWR _00252_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08908_ _04062_ _04065_ _04061_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__a21oi_1
X_09888_ _04734_ u_rf.reg7_q\[6\] _04722_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__mux2_1
X_08839_ _04007_ _04010_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_142_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ clknet_leaf_18_clk _00077_ net288 VGND VGND VPWR VPWR u_rf.reg0_q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_142_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10801_ _05248_ VGND VGND VPWR VPWR _00629_ sky130_fd_sc_hd__clkbuf_1
X_11781_ clknet_leaf_85_clk net164 net363 VGND VGND VPWR VPWR u_decod.pc0_q_i\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_323 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10732_ u_rf.reg18_q\[21\] _04983_ _05210_ VGND VGND VPWR VPWR _05212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ _05175_ VGND VGND VPWR VPWR _00564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12402_ clknet_leaf_40_clk _00439_ net278 VGND VGND VPWR VPWR u_rf.reg13_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10594_ u_rf.reg16_q\[20\] _04980_ _05138_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12333_ clknet_leaf_8_clk _00370_ net217 VGND VGND VPWR VPWR u_rf.reg11_q\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12264_ clknet_leaf_18_clk _00301_ net288 VGND VGND VPWR VPWR u_rf.reg9_q\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11215_ u_rf.reg25_q\[24\] _04989_ _05463_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__mux2_1
X_12195_ clknet_leaf_108_clk _00232_ net313 VGND VGND VPWR VPWR u_rf.reg7_q\[8\] sky130_fd_sc_hd__dfrtp_1
X_11146_ _05431_ VGND VGND VPWR VPWR _00791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11077_ _04770_ u_rf.reg23_q\[23\] _05391_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10028_ u_rf.reg8_q\[28\] _04486_ _04812_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11979_ clknet_leaf_75_clk net456 net368 VGND VGND VPWR VPWR u_decod.pc_q_o\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_737 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07170_ u_decod.rs2_data_q\[15\] _01289_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_601 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06121_ _01379_ _01383_ _01387_ _01391_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__or4b_2
XFILLER_0_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_120_clk clknet_4_3_0_clk VGND VGND VPWR VPWR clknet_leaf_120_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06052_ u_decod.rs1_data_q\[4\] u_decod.rs2_data_q\[4\] VGND VGND VPWR VPWR _01323_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_375 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout306 net307 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_4
Xfanout339 net340 VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_4
X_09811_ _04690_ VGND VGND VPWR VPWR _00197_ sky130_fd_sc_hd__clkbuf_1
Xfanout317 net318 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_2
Xfanout328 net330 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_4
X_09742_ _04653_ VGND VGND VPWR VPWR _00165_ sky130_fd_sc_hd__clkbuf_1
X_06954_ _02202_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[11\] sky130_fd_sc_hd__inv_2
X_05905_ u_decod.pc0_q_i\[31\] _01192_ _01195_ VGND VGND VPWR VPWR _01196_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09673_ _04615_ VGND VGND VPWR VPWR _00134_ sky130_fd_sc_hd__clkbuf_1
X_06885_ _01703_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__buf_2
X_08624_ u_rf.reg15_q\[21\] _03301_ _03303_ u_rf.reg24_q\[21\] _03806_ VGND VGND VPWR
+ VPWR _03807_ sky130_fd_sc_hd__a221o_1
X_05836_ _01098_ VGND VGND VPWR VPWR _01144_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ u_rf.reg4_q\[18\] _03224_ _03211_ u_rf.reg11_q\[18\] VGND VGND VPWR VPWR
+ _03741_ sky130_fd_sc_hd__a22o_1
X_05767_ _01068_ _01074_ VGND VGND VPWR VPWR _01090_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_38_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07506_ _02540_ _02732_ _01905_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08486_ u_rf.reg9_q\[15\] _03348_ _03349_ u_rf.reg20_q\[15\] VGND VGND VPWR VPWR
+ _03675_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07437_ u_rf.reg5_q\[20\] _02664_ _02665_ u_rf.reg19_q\[20\] _02666_ VGND VGND VPWR
+ VPWR _02667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07368_ u_rf.reg23_q\[19\] _01613_ _01609_ u_rf.reg12_q\[19\] _02599_ VGND VGND VPWR
+ VPWR _02600_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_264 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09107_ _04241_ _04236_ _04231_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06319_ u_rf.reg25_q\[0\] _01576_ _01581_ u_rf.reg30_q\[0\] _01588_ VGND VGND VPWR
+ VPWR _01589_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07299_ _01381_ _01400_ _02443_ _01387_ _01401_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_111_clk clknet_4_9_0_clk VGND VGND VPWR VPWR clknet_leaf_111_clk sky130_fd_sc_hd__clkbuf_16
X_09038_ _01366_ _01370_ _01383_ _01387_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__nand4_1
XFILLER_0_130_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11000_ u_rf.reg22_q\[19\] _04978_ _05344_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ clknet_leaf_71_clk _00988_ net354 VGND VGND VPWR VPWR u_rf.reg30_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_234 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12882_ clknet_leaf_41_clk _00919_ net298 VGND VGND VPWR VPWR u_rf.reg28_q\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_11902_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[23\] net347 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ clknet_leaf_112_clk net21 net321 VGND VGND VPWR VPWR u_decod.dec0.funct7\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_114_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11764_ clknet_leaf_66_clk _00056_ net349 VGND VGND VPWR VPWR u_rf.reg1_q\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_473 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11695_ _05722_ VGND VGND VPWR VPWR _01049_ sky130_fd_sc_hd__clkbuf_1
X_10715_ u_rf.reg18_q\[13\] _04966_ _05199_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10646_ _05166_ VGND VGND VPWR VPWR _00556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer5 _04028_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_212 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10577_ u_rf.reg16_q\[12\] _04964_ _05127_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_102_clk clknet_4_8_0_clk VGND VGND VPWR VPWR clknet_leaf_102_clk sky130_fd_sc_hd__clkbuf_16
X_12316_ clknet_leaf_128_clk _00353_ net236 VGND VGND VPWR VPWR u_rf.reg11_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12247_ clknet_leaf_50_clk _00284_ net308 VGND VGND VPWR VPWR u_rf.reg8_q\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ clknet_leaf_46_clk _00215_ net278 VGND VGND VPWR VPWR u_rf.reg6_q\[23\] sky130_fd_sc_hd__dfrtp_1
X_11129_ _05422_ VGND VGND VPWR VPWR _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06670_ u_rf.reg1_q\[5\] _01586_ _01635_ u_rf.reg9_q\[5\] VGND VGND VPWR VPWR _01930_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08340_ u_rf.reg6_q\[8\] _03387_ _03388_ u_rf.reg13_q\[8\] VGND VGND VPWR VPWR _03536_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_501 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08271_ u_rf.reg4_q\[5\] _03356_ _03311_ u_rf.reg1_q\[5\] _03469_ VGND VGND VPWR
+ VPWR _03470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07222_ u_decod.pc_q_o\[15\] u_decod.pc_q_o\[16\] _02335_ VGND VGND VPWR VPWR _02461_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_13_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_702 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07153_ _02225_ _02227_ _02278_ _02328_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__and4b_1
XFILLER_0_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_589 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06104_ _01362_ _01366_ _01370_ _01374_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__or4_1
XFILLER_0_14_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07084_ _02305_ _02306_ _02327_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06035_ u_decod.rs2_data_q\[9\] u_decod.rs1_data_q\[9\] VGND VGND VPWR VPWR _01306_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_126_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07986_ _01532_ u_decod.dec0.instr_i\[17\] _03170_ u_decod.rf_ff_rd_adr_q_i\[4\]
+ VGND VGND VPWR VPWR _03192_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_126_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _04642_ VGND VGND VPWR VPWR _00159_ sky130_fd_sc_hd__clkbuf_1
X_06937_ _01059_ _02183_ _02184_ _02185_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__o2bb2a_1
X_09656_ _04605_ VGND VGND VPWR VPWR _00127_ sky130_fd_sc_hd__clkbuf_1
X_08607_ _03784_ _03786_ _03788_ _03790_ VGND VGND VPWR VPWR _03791_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_2_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ _02113_ _02115_ _02117_ _02119_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__or4_1
XFILLER_0_139_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05819_ _01129_ _01106_ _01130_ VGND VGND VPWR VPWR _01131_ sky130_fd_sc_hd__and3b_1
X_09587_ u_decod.rf_ff_rd_adr_q_i\[0\] _04424_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand2_2
X_06799_ u_decod.pc_q_o\[6\] u_decod.pc_q_o\[7\] u_decod.pc_q_o\[8\] _01917_ VGND
+ VGND VPWR VPWR _02054_ sky130_fd_sc_hd__and4_2
X_08538_ u_rf.reg0_q\[17\] _03175_ _03328_ u_rf.reg12_q\[17\] _03724_ VGND VGND VPWR
+ VPWR _03725_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08469_ u_rf.reg16_q\[14\] _03248_ _03249_ u_rf.reg5_q\[14\] VGND VGND VPWR VPWR
+ _03659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10500_ _04740_ u_rf.reg15_q\[9\] _05078_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11480_ _05608_ VGND VGND VPWR VPWR _00948_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_521 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10431_ _05051_ VGND VGND VPWR VPWR _00456_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10362_ _04738_ u_rf.reg13_q\[8\] _05006_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__mux2_1
X_10293_ u_rf.reg12_q\[15\] _04970_ _04960_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__mux2_1
X_12101_ clknet_leaf_125_clk _00138_ net239 VGND VGND VPWR VPWR u_rf.reg4_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12032_ clknet_leaf_114_clk u_decod.exe_ff_res_data_i\[12\] net330 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12934_ clknet_leaf_138_clk _00971_ net210 VGND VGND VPWR VPWR u_rf.reg30_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12865_ clknet_leaf_117_clk _00902_ net325 VGND VGND VPWR VPWR u_rf.reg28_q\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11816_ clknet_leaf_98_clk net3 net331 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_12796_ clknet_leaf_126_clk _00833_ net240 VGND VGND VPWR VPWR u_rf.reg26_q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11747_ clknet_leaf_130_clk _00039_ net234 VGND VGND VPWR VPWR u_rf.reg1_q\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11678_ _05713_ VGND VGND VPWR VPWR _01041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_318 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10629_ _05157_ VGND VGND VPWR VPWR _00548_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_362 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07840_ _03014_ _03052_ _01481_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__mux2_1
X_07771_ u_rf.reg1_q\[27\] _02604_ _02367_ u_rf.reg14_q\[27\] VGND VGND VPWR VPWR
+ _02987_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_108_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09510_ u_rf.reg1_q\[28\] _04486_ _04518_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06722_ u_rf.reg19_q\[6\] _01593_ _01644_ u_rf.reg20_q\[6\] VGND VGND VPWR VPWR _01980_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09441_ u_rf.reg2_q\[29\] _04488_ _04470_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_121_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06653_ net37 _01489_ _01490_ net54 VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__a22o_1
X_09372_ u_decod.rf_ff_res_data_i\[7\] VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__buf_2
X_06584_ u_rf.reg9_q\[3\] _01635_ _01656_ u_rf.reg10_q\[3\] VGND VGND VPWR VPWR _01848_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08323_ _03512_ _03514_ _03517_ _03519_ VGND VGND VPWR VPWR _03520_ sky130_fd_sc_hd__or4_1
XFILLER_0_145_821 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_865 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08254_ u_rf.reg0_q\[4\] _03176_ _03329_ u_rf.reg12_q\[4\] _03453_ VGND VGND VPWR
+ VPWR _03454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_729 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07205_ net99 net39 _01064_ _01067_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__and4_1
X_08185_ _03304_ VGND VGND VPWR VPWR _03387_ sky130_fd_sc_hd__buf_6
XFILLER_0_132_559 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07136_ u_rf.reg11_q\[14\] _02375_ _02376_ u_rf.reg13_q\[14\] _02377_ VGND VGND VPWR
+ VPWR _02378_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07067_ u_rf.reg15_q\[13\] _01601_ _01608_ u_rf.reg12_q\[13\] _02310_ VGND VGND VPWR
+ VPWR _02311_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06018_ u_decod.rs1_data_q\[15\] VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09708_ u_rf.reg4_q\[23\] _04476_ _04630_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__mux2_1
X_07969_ _03174_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__buf_6
X_10980_ _05343_ VGND VGND VPWR VPWR _00713_ sky130_fd_sc_hd__clkbuf_1
X_09639_ u_rf.reg3_q\[23\] _04476_ _04593_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12650_ clknet_leaf_29_clk _00687_ net260 VGND VGND VPWR VPWR u_rf.reg21_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_629 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _05672_ VGND VGND VPWR VPWR _01005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_681 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12581_ clknet_leaf_124_clk _00618_ net239 VGND VGND VPWR VPWR u_rf.reg19_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_854 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11532_ _04749_ u_rf.reg30_q\[13\] _05632_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11463_ _05599_ VGND VGND VPWR VPWR _00940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10414_ _04719_ u_rf.reg14_q\[0\] _05042_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11394_ u_rf.reg28_q\[12\] u_decod.rf_ff_res_data_i\[12\] _05560_ VGND VGND VPWR
+ VPWR _05563_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10345_ _05005_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__buf_8
XFILLER_0_21_579 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10276_ u_decod.rf_ff_res_data_i\[10\] VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__buf_2
X_12015_ clknet_leaf_76_clk u_exe.bu_pc_res\[28\] net368 VGND VGND VPWR VPWR u_exe.pc_data_q\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12917_ clknet_leaf_47_clk _00954_ net301 VGND VGND VPWR VPWR u_rf.reg29_q\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12848_ clknet_leaf_31_clk _00885_ net264 VGND VGND VPWR VPWR u_rf.reg27_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12779_ clknet_leaf_2_clk _00816_ net223 VGND VGND VPWR VPWR u_rf.reg25_q\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_813 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_822 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09990_ _04789_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__buf_6
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08941_ _01380_ u_decod.branch_imm_q_o\[17\] _04097_ VGND VGND VPWR VPWR _04098_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08872_ u_decod.rs1_data_q\[6\] u_decod.branch_imm_q_o\[6\] _04038_ _04031_ VGND
+ VGND VPWR VPWR _04039_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_4_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07823_ u_rf.reg18_q\[28\] _01787_ _02367_ u_rf.reg14_q\[28\] _03036_ VGND VGND VPWR
+ VPWR _03037_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07754_ _01485_ _02957_ _02958_ _02970_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07685_ u_decod.rf_ff_res_data_i\[25\] _01550_ _02743_ _02884_ _02904_ VGND VGND
+ VPWR VPWR _02905_ sky130_fd_sc_hd__a221o_1
X_06705_ _01484_ _01962_ _01963_ _01428_ _01329_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__a32o_1
XFILLER_0_149_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09424_ _04477_ VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_91_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_06636_ _01802_ _01853_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06567_ u_decod.dec0.instr_i\[10\] _01226_ _01715_ u_decod.dec0.instr_i\[23\] VGND
+ VGND VPWR VPWR _01831_ sky130_fd_sc_hd__a22o_1
X_09355_ u_rf.reg2_q\[1\] _04430_ _04428_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_785 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06498_ u_decod.instr_operation_q\[0\] _01259_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__nand2_4
X_08306_ u_rf.reg18_q\[7\] _03353_ _03355_ u_rf.reg23_q\[7\] _03502_ VGND VGND VPWR
+ VPWR _03503_ sky130_fd_sc_hd__a221o_1
X_09286_ _04385_ u_decod.rs2_data_q\[6\] _04386_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08237_ u_rf.reg22_q\[4\] _03275_ _03277_ u_rf.reg3_q\[4\] VGND VGND VPWR VPWR _03437_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08168_ u_rf.reg1_q\[1\] _03310_ _03312_ u_rf.reg14_q\[1\] VGND VGND VPWR VPWR _03371_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08099_ _03302_ VGND VGND VPWR VPWR _03303_ sky130_fd_sc_hd__buf_8
X_07119_ u_rf.reg19_q\[14\] _01595_ _01650_ u_rf.reg4_q\[14\] VGND VGND VPWR VPWR
+ _02361_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_765 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10130_ u_rf.reg10_q\[11\] _04451_ _04874_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10061_ _04839_ VGND VGND VPWR VPWR _00298_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10963_ u_rf.reg22_q\[1\] _04941_ _05333_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_82_clk clknet_4_14_0_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12702_ clknet_leaf_123_clk _00739_ net232 VGND VGND VPWR VPWR u_rf.reg23_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10894_ _05298_ VGND VGND VPWR VPWR _00672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12633_ clknet_leaf_62_clk _00670_ net342 VGND VGND VPWR VPWR u_rf.reg20_q\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12564_ clknet_leaf_24_clk _00601_ net267 VGND VGND VPWR VPWR u_rf.reg18_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11515_ _04732_ u_rf.reg30_q\[5\] _05621_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__mux2_1
X_12495_ clknet_leaf_38_clk _00532_ net274 VGND VGND VPWR VPWR u_rf.reg16_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11446_ _05590_ VGND VGND VPWR VPWR _00932_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_237 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11377_ u_rf.reg28_q\[4\] net512 _05549_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__mux2_1
X_10328_ _04994_ VGND VGND VPWR VPWR _00410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10259_ u_rf.reg12_q\[4\] _04947_ _04939_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_clk clknet_4_15_0_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07470_ u_rf.reg30_q\[21\] _01581_ _02419_ u_rf.reg28_q\[21\] VGND VGND VPWR VPWR
+ _02698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06421_ _01474_ _01452_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09140_ _04268_ _04269_ VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06352_ _01621_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__buf_6
XFILLER_0_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09071_ u_decod.pc_q_o\[2\] u_decod.branch_imm_q_o\[2\] VGND VGND VPWR VPWR _04211_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06283_ u_decod.dec0.instr_i\[20\] _01552_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__nor2_2
XFILLER_0_114_312 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08022_ _03208_ _03215_ _03221_ _03227_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__or4_1
XFILLER_0_72_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_576 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09973_ _04792_ VGND VGND VPWR VPWR _00257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08924_ _04042_ _04083_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__nor2_1
XFILLER_0_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08855_ u_decod.rs1_data_q\[6\] u_decod.branch_imm_q_o\[6\] VGND VGND VPWR VPWR _04024_
+ sky130_fd_sc_hd__and2_1
X_08786_ u_rf.reg0_q\[29\] _03175_ _03357_ u_rf.reg17_q\[29\] _03960_ VGND VGND VPWR
+ VPWR _03961_ sky130_fd_sc_hd__a221o_1
X_07806_ u_decod.dec0.funct7\[3\] _01224_ _02646_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _02952_ _02954_ VGND VGND VPWR VPWR u_decod.rs2_data_nxt\[26\] sky130_fd_sc_hd__xnor2_1
X_05998_ u_decod.rs2_data_q\[31\] _01267_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_64_clk clknet_4_12_0_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_354 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_905 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07668_ u_rf.reg1_q\[25\] _01586_ _01671_ u_rf.reg27_q\[25\] _02887_ VGND VGND VPWR
+ VPWR _02888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07599_ _01357_ _01393_ _01407_ _01280_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__a211o_1
X_09407_ u_rf.reg2_q\[18\] _04465_ _04449_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06619_ u_rf.reg14_q\[4\] _01658_ _01670_ u_rf.reg27_q\[4\] VGND VGND VPWR VPWR _01881_
+ sky130_fd_sc_hd__a22o_1
X_09338_ _04409_ u_decod.rs2_data_q\[30\] _04410_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__and3_1
XFILLER_0_75_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_301 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09269_ _04373_ _04379_ _04378_ _04377_ VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_106_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11300_ _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_893 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12280_ clknet_leaf_53_clk _00317_ net302 VGND VGND VPWR VPWR u_rf.reg9_q\[29\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11231_ _04682_ _04825_ _05295_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__and3_2
XFILLER_0_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11162_ _05439_ VGND VGND VPWR VPWR _00799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10113_ u_rf.reg10_q\[3\] _04434_ _04863_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__mux2_1
X_11093_ _04786_ u_rf.reg23_q\[31\] _05368_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__mux2_1
X_10044_ _04830_ VGND VGND VPWR VPWR _00290_ sky130_fd_sc_hd__clkbuf_1
Xhold61 u_decod.pc0_q_i\[30\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 u_decod.dec0.funct7\[1\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 u_decod.exe_ff_rd_adr_q_i\[3\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold94 u_exe.pc_data_q\[10\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_55_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
X_11995_ clknet_leaf_85_clk u_exe.bu_pc_res\[8\] net363 VGND VGND VPWR VPWR u_exe.pc_data_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10946_ _05325_ VGND VGND VPWR VPWR _00697_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_404 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10877_ _05288_ VGND VGND VPWR VPWR _00665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_757 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12616_ clknet_leaf_21_clk _00653_ net282 VGND VGND VPWR VPWR u_rf.reg20_q\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_891 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_632 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12547_ clknet_leaf_105_clk _00584_ net319 VGND VGND VPWR VPWR u_rf.reg18_q\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_3 _01206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12478_ clknet_leaf_134_clk _00515_ net232 VGND VGND VPWR VPWR u_rf.reg16_q\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_427 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11429_ u_rf.reg28_q\[29\] u_decod.rf_ff_res_data_i\[29\] _05571_ VGND VGND VPWR
+ VPWR _05581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_315 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06970_ u_rf.reg17_q\[11\] _01630_ _01635_ u_rf.reg9_q\[11\] VGND VGND VPWR VPWR
+ _02218_ sky130_fd_sc_hd__a22o_1
X_05921_ u_decod.dec0.funct3\[1\] u_decod.dec0.funct3\[2\] _01209_ _01210_ VGND VGND
+ VPWR VPWR _01211_ sky130_fd_sc_hd__or4_1
X_05852_ u_decod.pc0_q_i\[18\] _01153_ VGND VGND VPWR VPWR _01156_ sky130_fd_sc_hd__or2_1
X_08640_ u_rf.reg7_q\[22\] _03369_ _03313_ u_rf.reg14_q\[22\] _03821_ VGND VGND VPWR
+ VPWR _03822_ sky130_fd_sc_hd__a221o_1
Xrebuffer26 net401 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer15 u_decod.pc0_q_i\[3\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_4_7_0_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
Xrebuffer37 _01129_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__dlygate4sd1_1
X_05783_ net441 _01099_ _01101_ net76 _01103_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__a221o_2
X_08571_ u_rf.reg4_q\[19\] _03356_ _03357_ u_rf.reg17_q\[19\] _03755_ VGND VGND VPWR
+ VPWR _03756_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_505 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07522_ u_rf.reg6_q\[22\] _01557_ _02604_ u_rf.reg1_q\[22\] _02747_ VGND VGND VPWR
+ VPWR _02748_ sky130_fd_sc_hd__a221o_1
X_07453_ _02580_ _02680_ _02681_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__mux2_1
X_06404_ _01673_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09123_ _04047_ _04207_ _04208_ _04255_ VGND VGND VPWR VPWR u_exe.bu_pc_res\[9\]
+ sky130_fd_sc_hd__a2bb2o_1
X_07384_ _01772_ u_decod.exe_ff_res_data_i\[19\] _02615_ VGND VGND VPWR VPWR _02616_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_755 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_643 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_552 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06335_ _01604_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__buf_8
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ _04195_ VGND VGND VPWR VPWR _04196_ sky130_fd_sc_hd__buf_2
X_06266_ u_decod.rf_ff_rd_adr_q_i\[3\] VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08005_ _03171_ _03201_ _03209_ VGND VGND VPWR VPWR _03211_ sky130_fd_sc_hd__and3_4
XFILLER_0_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06197_ _01467_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_696 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_493 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09956_ _04780_ u_rf.reg7_q\[28\] _04764_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ _04067_ _04068_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nor2_1
X_09887_ u_decod.rf_ff_res_data_i\[6\] VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__buf_2
X_08838_ _04008_ _04009_ VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08769_ u_rf.reg6_q\[28\] _03304_ _03306_ u_rf.reg13_q\[28\] VGND VGND VPWR VPWR
+ _03945_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_142_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_5_0_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10800_ u_rf.reg19_q\[21\] _04983_ _05246_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__mux2_1
X_11780_ clknet_leaf_85_clk net163 net363 VGND VGND VPWR VPWR u_decod.pc0_q_i\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_713 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10731_ _05211_ VGND VGND VPWR VPWR _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10662_ u_rf.reg17_q\[20\] _04980_ _05174_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__mux2_1
X_12401_ clknet_leaf_53_clk _00438_ net302 VGND VGND VPWR VPWR u_rf.reg13_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10593_ _05115_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_11_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_766 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12332_ clknet_leaf_14_clk _00369_ net246 VGND VGND VPWR VPWR u_rf.reg11_q\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_224 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12263_ clknet_leaf_4_clk _00300_ net212 VGND VGND VPWR VPWR u_rf.reg9_q\[12\] sky130_fd_sc_hd__dfrtp_1
X_11214_ _05467_ VGND VGND VPWR VPWR _00823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12194_ clknet_leaf_129_clk _00231_ net235 VGND VGND VPWR VPWR u_rf.reg7_q\[7\] sky130_fd_sc_hd__dfrtp_1
X_11145_ u_rf.reg24_q\[23\] _04987_ _05427_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__mux2_1
X_11076_ _05394_ VGND VGND VPWR VPWR _00758_ sky130_fd_sc_hd__clkbuf_1
X_10027_ _04820_ VGND VGND VPWR VPWR _00283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_4_4_0_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11978_ clknet_leaf_73_clk net452 net369 VGND VGND VPWR VPWR u_decod.pc_q_o\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_19_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10929_ _05316_ VGND VGND VPWR VPWR _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06120_ _01389_ _01390_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__nor2_2
XFILLER_0_152_793 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06051_ u_decod.rs1_data_q\[4\] u_decod.rs2_data_q\[4\] VGND VGND VPWR VPWR _01322_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_41_246 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_281 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_145 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout307 net309 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__buf_2
XFILLER_0_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09810_ u_rf.reg6_q\[5\] _04438_ _04684_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__mux2_1
Xfanout329 net330 VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_4
Xfanout318 net334 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__buf_2
XFILLER_0_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09741_ u_rf.reg5_q\[5\] _04438_ _04647_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__mux2_1
X_06953_ _01437_ _02181_ _02187_ _02201_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_05904_ u_decod.pc0_q_i\[31\] _01192_ _01106_ VGND VGND VPWR VPWR _01195_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09672_ u_rf.reg4_q\[6\] _04440_ _04608_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__mux2_1
X_06884_ _01345_ _01305_ _01308_ _01341_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__or4_1
X_08623_ u_rf.reg6_q\[21\] _03305_ _03307_ u_rf.reg13_q\[21\] VGND VGND VPWR VPWR
+ _03806_ sky130_fd_sc_hd__a22o_1
X_05835_ u_decod.pc0_q_i\[14\] _01139_ VGND VGND VPWR VPWR _01143_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_clk clknet_4_6_0_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_124_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08554_ _03733_ _03735_ _03737_ _03739_ VGND VGND VPWR VPWR _03740_ sky130_fd_sc_hd__or4_1
XFILLER_0_11_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05766_ _01085_ _01088_ VGND VGND VPWR VPWR _01089_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_38_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_644 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07505_ _01371_ _01292_ u_decod.rs1_data_q\[6\] _01747_ _01467_ _01461_ VGND VGND
+ VPWR VPWR _02732_ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08485_ u_rf.reg18_q\[15\] _03353_ _03355_ u_rf.reg23_q\[15\] _03673_ VGND VGND VPWR
+ VPWR _03674_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07436_ u_rf.reg16_q\[20\] _01565_ _01631_ u_rf.reg17_q\[20\] VGND VGND VPWR VPWR
+ _02666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_738 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07367_ u_rf.reg16_q\[19\] _01564_ _01670_ u_rf.reg27_q\[19\] VGND VGND VPWR VPWR
+ _02599_ sky130_fd_sc_hd__a22o_1
X_09106_ _04233_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_06318_ u_rf.reg11_q\[0\] _01584_ _01587_ u_rf.reg1_q\[0\] VGND VGND VPWR VPWR _01588_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09037_ _01355_ _01352_ _02588_ _01391_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__or4_1
X_07298_ _01387_ _02532_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_657 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06249_ u_decod.dec0.instr_i\[23\] u_decod.exe_ff_rd_adr_q_i\[3\] VGND VGND VPWR
+ VPWR _01519_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_144_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_09939_ _04769_ VGND VGND VPWR VPWR _00246_ sky130_fd_sc_hd__clkbuf_1
X_12950_ clknet_leaf_50_clk _00987_ net309 VGND VGND VPWR VPWR u_rf.reg30_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_12881_ clknet_leaf_53_clk _00918_ net302 VGND VGND VPWR VPWR u_rf.reg28_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11901_ clknet_leaf_90_clk u_decod.rs2_data_nxt\[22\] net345 VGND VGND VPWR VPWR
+ u_decod.rs2_data_q\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ clknet_leaf_112_clk net20 net321 VGND VGND VPWR VPWR u_decod.dec0.funct7\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_11763_ clknet_leaf_39_clk _00055_ net277 VGND VGND VPWR VPWR u_rf.reg1_q\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11694_ u_decod.branch_imm_q_o\[25\] _02884_ _05717_ VGND VGND VPWR VPWR _05722_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10714_ _05202_ VGND VGND VPWR VPWR _00588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10645_ u_rf.reg17_q\[12\] _04964_ _05163_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer6 net379 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12315_ clknet_leaf_12_clk _00352_ net242 VGND VGND VPWR VPWR u_rf.reg11_q\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10576_ _05129_ VGND VGND VPWR VPWR _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_268 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12246_ clknet_leaf_50_clk _00283_ net308 VGND VGND VPWR VPWR u_rf.reg8_q\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_139_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12177_ clknet_leaf_56_clk _00214_ net293 VGND VGND VPWR VPWR u_rf.reg6_q\[22\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_75_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11128_ u_rf.reg24_q\[15\] _04970_ _05416_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11059_ _05385_ VGND VGND VPWR VPWR _00750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_13 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08270_ u_rf.reg31_q\[5\] _03210_ _03343_ u_rf.reg26_q\[5\] VGND VGND VPWR VPWR _03469_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07221_ _01505_ _02451_ _02453_ _02459_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__a211o_1
X_07152_ _02357_ u_decod.exe_ff_res_data_i\[14\] _02393_ VGND VGND VPWR VPWR _02394_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_714 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06103_ _01372_ _01373_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07083_ u_decod.rf_ff_res_data_i\[13\] _01549_ u_decod.exe_ff_res_data_i\[13\] _01713_
+ _02326_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_8_clk clknet_4_1_0_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
X_06034_ u_decod.rs2_data_q\[9\] u_decod.rs1_data_q\[9\] VGND VGND VPWR VPWR _01305_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07985_ u_decod.dec0.instr_i\[18\] VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_126_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09724_ u_rf.reg4_q\[31\] _04492_ _04607_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__mux2_1
X_06936_ u_decod.pc_q_o\[9\] u_decod.pc_q_o\[10\] u_decod.pc_q_o\[11\] _02054_ VGND
+ VGND VPWR VPWR _02185_ sky130_fd_sc_hd__and4_2
X_09655_ u_rf.reg3_q\[31\] _04492_ _04570_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__mux2_1
X_06867_ u_rf.reg12_q\[9\] _01607_ _01672_ u_rf.reg2_q\[9\] _02118_ VGND VGND VPWR
+ VPWR _02119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08606_ u_rf.reg0_q\[20\] _03420_ _03421_ u_rf.reg12_q\[20\] _03789_ VGND VGND VPWR
+ VPWR _03790_ sky130_fd_sc_hd__a221o_1
X_05818_ u_decod.pc0_q_i\[9\] net385 u_decod.pc0_q_i\[10\] VGND VGND VPWR VPWR _01130_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _04567_ VGND VGND VPWR VPWR _00095_ sky130_fd_sc_hd__clkbuf_1
X_06798_ u_decod.pc_q_o\[8\] _02006_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08537_ u_rf.reg28_q\[17\] _03242_ _03243_ u_rf.reg2_q\[17\] VGND VGND VPWR VPWR
+ _03724_ sky130_fd_sc_hd__a22o_1
X_05749_ u_decod.dec0.instr_i\[3\] VGND VGND VPWR VPWR _01072_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08468_ u_rf.reg0_q\[14\] _03175_ _03328_ u_rf.reg12_q\[14\] _03657_ VGND VGND VPWR
+ VPWR _03658_ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_07419_ u_rf.reg13_q\[20\] _01598_ _01592_ u_rf.reg18_q\[20\] _02648_ VGND VGND VPWR
+ VPWR _02649_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10430_ _04738_ u_rf.reg14_q\[8\] _05042_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__mux2_1
X_08399_ u_rf.reg31_q\[11\] _03504_ _03505_ u_rf.reg11_q\[11\] _03591_ VGND VGND VPWR
+ VPWR _03592_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_154_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _05014_ VGND VGND VPWR VPWR _00423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10292_ u_decod.rf_ff_res_data_i\[15\] VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12100_ clknet_leaf_107_clk _00137_ net314 VGND VGND VPWR VPWR u_rf.reg4_q\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_57_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12031_ clknet_leaf_114_clk u_decod.exe_ff_res_data_i\[11\] net328 VGND VGND VPWR
+ VPWR u_decod.rf_ff_res_data_i\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ clknet_leaf_120_clk _00970_ net249 VGND VGND VPWR VPWR u_rf.reg30_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12864_ clknet_leaf_114_clk _00901_ net327 VGND VGND VPWR VPWR u_rf.reg28_q\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_157_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_841 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11815_ clknet_leaf_114_clk net2 net328 VGND VGND VPWR VPWR u_decod.dec0.instr_i\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12795_ clknet_leaf_122_clk _00832_ net248 VGND VGND VPWR VPWR u_rf.reg26_q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11746_ clknet_leaf_119_clk _00038_ net251 VGND VGND VPWR VPWR u_rf.reg1_q\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11677_ u_decod.branch_imm_q_o\[17\] _02509_ _05696_ VGND VGND VPWR VPWR _05713_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10628_ u_rf.reg17_q\[4\] _04947_ _05152_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_47_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10559_ _05120_ VGND VGND VPWR VPWR _00515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12229_ clknet_leaf_125_clk _00266_ net239 VGND VGND VPWR VPWR u_rf.reg8_q\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_07770_ u_rf.reg0_q\[27\] _01664_ _02371_ u_rf.reg15_q\[27\] _02985_ VGND VGND VPWR
+ VPWR _02986_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06721_ u_rf.reg13_q\[6\] _01597_ _01600_ u_rf.reg15_q\[6\] _01978_ VGND VGND VPWR
+ VPWR _01979_ sky130_fd_sc_hd__a221o_1
X_09440_ u_decod.rf_ff_res_data_i\[29\] VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_56_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06652_ _01423_ _01870_ _01912_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__o21ai_1
X_09371_ _04441_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06583_ u_rf.reg0_q\[3\] _01663_ _01645_ u_rf.reg20_q\[3\] _01846_ VGND VGND VPWR
+ VPWR _01847_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08322_ u_rf.reg0_q\[7\] _03176_ _03329_ u_rf.reg12_q\[7\] _03518_ VGND VGND VPWR
+ VPWR _03519_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08253_ u_rf.reg28_q\[4\] _03331_ _03333_ u_rf.reg2_q\[4\] VGND VGND VPWR VPWR _03453_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07204_ _01290_ _01294_ _01356_ _01391_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_74_477 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_365 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08184_ u_rf.reg7_q\[2\] _03314_ _03315_ u_rf.reg25_q\[2\] _03385_ VGND VGND VPWR
+ VPWR _03386_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_65_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07135_ u_rf.reg30_q\[14\] _01580_ _01592_ u_rf.reg18_q\[14\] VGND VGND VPWR VPWR
+ _02377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07066_ u_rf.reg25_q\[13\] _01575_ _01624_ u_rf.reg28_q\[13\] VGND VGND VPWR VPWR
+ _02310_ sky130_fd_sc_hd__a22o_1
X_06017_ _01274_ _01287_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07968_ _03171_ _03172_ _03173_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__and3_4
X_09707_ _04633_ VGND VGND VPWR VPWR _00150_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_74_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_06919_ u_rf.reg29_q\[10\] _01626_ _01637_ u_rf.reg21_q\[10\] _02168_ VGND VGND VPWR
+ VPWR _02169_ sky130_fd_sc_hd__a221o_1
X_07899_ u_rf.reg1_q\[30\] _02604_ _02419_ u_rf.reg28_q\[30\] _03108_ VGND VGND VPWR
+ VPWR _03109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09638_ _04596_ VGND VGND VPWR VPWR _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ u_rf.reg0_q\[23\] _04476_ _04555_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _04749_ u_rf.reg31_q\[13\] _05668_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_411 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ clknet_leaf_111_clk _00617_ net316 VGND VGND VPWR VPWR u_rf.reg19_q\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11531_ _05635_ VGND VGND VPWR VPWR _00972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_83_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11462_ _04747_ u_rf.reg29_q\[12\] _05596_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10413_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_59_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11393_ _05562_ VGND VGND VPWR VPWR _00907_ sky130_fd_sc_hd__clkbuf_1
X_10344_ _01534_ _04424_ _04423_ _04936_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_72_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10275_ _04958_ VGND VGND VPWR VPWR _00393_ sky130_fd_sc_hd__clkbuf_1
X_12014_ clknet_leaf_76_clk u_exe.bu_pc_res\[27\] net369 VGND VGND VPWR VPWR u_exe.pc_data_q\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_92_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12916_ clknet_leaf_23_clk _00953_ net268 VGND VGND VPWR VPWR u_rf.reg29_q\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12847_ clknet_leaf_37_clk _00884_ net273 VGND VGND VPWR VPWR u_rf.reg27_q\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12778_ clknet_leaf_29_clk _00815_ net260 VGND VGND VPWR VPWR u_rf.reg25_q\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_809 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11729_ clknet_leaf_35_clk _00021_ net271 VGND VGND VPWR VPWR u_rf.reg2_q\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_825 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_869 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_398 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_834 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08940_ _01380_ u_decod.branch_imm_q_o\[17\] u_decod.branch_imm_q_o\[16\] _01388_
+ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08871_ u_decod.rs1_data_q\[7\] u_decod.branch_imm_q_o\[7\] VGND VGND VPWR VPWR _04038_
+ sky130_fd_sc_hd__or2_1
X_07822_ u_rf.reg16_q\[28\] _02307_ _01784_ u_rf.reg24_q\[28\] VGND VGND VPWR VPWR
+ _03036_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_4_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07753_ net133 _02959_ _02963_ _02969_ VGND VGND VPWR VPWR _02970_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07684_ _01680_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__and2_2
X_06704_ u_decod.pc_q_o\[6\] _01917_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__nand2_1
X_09423_ u_rf.reg2_q\[23\] _04476_ _04470_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__mux2_1
X_06635_ _01093_ _01090_ _01896_ _01079_ _01237_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__a221o_4
XFILLER_0_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09354_ u_decod.rf_ff_res_data_i\[1\] VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_06566_ _01830_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[3\] sky130_fd_sc_hd__buf_1
XFILLER_0_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08305_ u_rf.reg4_q\[7\] _03356_ _03357_ u_rf.reg17_q\[7\] VGND VGND VPWR VPWR _03502_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_641 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_701 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_530 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09285_ _04389_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__buf_1
X_06497_ u_decod.instr_unit_q\[2\] _01056_ VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__nand2_4
XFILLER_0_145_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08236_ u_rf.reg18_q\[4\] _03262_ _03263_ u_rf.reg23_q\[4\] _03435_ VGND VGND VPWR
+ VPWR _03436_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_134_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08167_ _03230_ VGND VGND VPWR VPWR _03370_ sky130_fd_sc_hd__buf_8
X_07118_ _01636_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__clkbuf_8
X_08098_ _03238_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_54_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_07049_ _01460_ _01903_ _02293_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10060_ u_rf.reg9_q\[10\] _04448_ _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_845 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10962_ _05334_ VGND VGND VPWR VPWR _00704_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12701_ clknet_leaf_14_clk _00738_ net246 VGND VGND VPWR VPWR u_rf.reg23_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10893_ u_rf.reg21_q\[0\] _04935_ _05297_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12632_ clknet_leaf_52_clk _00669_ net351 VGND VGND VPWR VPWR u_rf.reg20_q\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_449 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12563_ clknet_leaf_68_clk _00600_ net351 VGND VGND VPWR VPWR u_rf.reg18_q\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12494_ clknet_leaf_7_clk _00531_ net218 VGND VGND VPWR VPWR u_rf.reg16_q\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11514_ _05626_ VGND VGND VPWR VPWR _00964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11445_ _04730_ u_rf.reg29_q\[4\] _05585_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11376_ _05553_ VGND VGND VPWR VPWR _00899_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10327_ u_rf.reg12_q\[26\] _04993_ _04981_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10258_ u_decod.rf_ff_res_data_i\[4\] VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__buf_2
X_10189_ _04907_ VGND VGND VPWR VPWR _00358_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_85_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_46 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06420_ _01465_ _01687_ _01688_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_06351_ _01620_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__buf_8
XFILLER_0_154_460 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_803 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09070_ u_decod.pc_q_o\[2\] u_decod.branch_imm_q_o\[2\] VGND VGND VPWR VPWR _04210_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06282_ u_decod.dec0.instr_i\[21\] VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__inv_2
XFILLER_0_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08021_ u_rf.reg18_q\[31\] _03222_ _03223_ u_rf.reg23_q\[31\] _03226_ VGND VGND VPWR
+ VPWR _03227_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_116_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_880 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09972_ u_rf.reg8_q\[1\] _04430_ _04790_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08923_ _04081_ _04082_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08854_ u_decod.rs1_data_q\[6\] u_decod.branch_imm_q_o\[6\] VGND VGND VPWR VPWR _04023_
+ sky130_fd_sc_hd__nor2_1
X_08785_ u_rf.reg31_q\[29\] _03289_ _03332_ u_rf.reg2_q\[29\] VGND VGND VPWR VPWR
+ _03960_ sky130_fd_sc_hd__a22o_1
X_07805_ _03019_ VGND VGND VPWR VPWR u_decod.exe_ff_res_data_i\[28\] sky130_fd_sc_hd__inv_2
X_05997_ u_decod.rs2_data_q\[31\] _01267_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__and2_1
X_07736_ _02864_ _02953_ net200 VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_366 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_07667_ u_rf.reg7_q\[25\] _01560_ _01644_ u_rf.reg20_q\[25\] VGND VGND VPWR VPWR
+ _02887_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07598_ _02818_ _01375_ _02635_ _02819_ _02820_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__a221o_1
X_09406_ u_decod.rf_ff_res_data_i\[18\] VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06618_ u_rf.reg12_q\[4\] _01608_ _01673_ u_rf.reg2_q\[4\] _01879_ VGND VGND VPWR
+ VPWR _01880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09337_ _04417_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__buf_1
X_06549_ _01811_ _01813_ _01765_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09268_ _04377_ _04378_ _04379_ _04373_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08219_ _03175_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__buf_8
XFILLER_0_7_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09199_ _04307_ _04314_ _04312_ _04311_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11230_ _05475_ VGND VGND VPWR VPWR _00831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11161_ u_rf.reg24_q\[31\] _05003_ _05404_ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10112_ _04866_ VGND VGND VPWR VPWR _00322_ sky130_fd_sc_hd__clkbuf_1
X_11092_ _05402_ VGND VGND VPWR VPWR _00766_ sky130_fd_sc_hd__clkbuf_1
X_10043_ u_rf.reg9_q\[2\] _04432_ _04827_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__mux2_1
Xhold62 u_decod.pc0_q_i\[31\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_1
Xhold73 u_decod.exe_ff_rd_adr_q_i\[0\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 u_decod.pc0_q_i\[18\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold84 u_decod.dec0.funct7\[0\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ clknet_leaf_85_clk u_exe.bu_pc_res\[7\] net363 VGND VGND VPWR VPWR u_exe.pc_data_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ u_rf.reg21_q\[25\] _04991_ _05319_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_11_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_725 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10876_ u_rf.reg20_q\[25\] _04991_ _05282_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_769 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12615_ clknet_leaf_5_clk _00652_ net214 VGND VGND VPWR VPWR u_rf.reg20_q\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_685 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12546_ clknet_leaf_130_clk _00583_ net230 VGND VGND VPWR VPWR u_rf.reg18_q\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12477_ clknet_leaf_14_clk _00514_ net244 VGND VGND VPWR VPWR u_rf.reg16_q\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11428_ _05580_ VGND VGND VPWR VPWR _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_4 _01469_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11359_ _04780_ u_rf.reg27_q\[28\] _05535_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_837 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ u_decod.dec0.funct3\[0\] u_decod.dec0.funct7\[6\] u_decod.dec0.instr_i\[20\]
+ VGND VGND VPWR VPWR _01210_ sky130_fd_sc_hd__or3_1
X_05851_ net501 _01142_ _01132_ net73 _01155_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__a221o_1
Xrebuffer27 net402 VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
Xrebuffer16 u_decod.pc0_q_i\[2\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__buf_1
X_08570_ u_rf.reg18_q\[19\] _03352_ _03354_ u_rf.reg23_q\[19\] VGND VGND VPWR VPWR
+ _03755_ sky130_fd_sc_hd__a22o_1
X_07521_ u_rf.reg25_q\[22\] _01576_ _02368_ u_rf.reg26_q\[22\] VGND VGND VPWR VPWR
+ _02747_ sky130_fd_sc_hd__a22o_1
X_05782_ u_decod.flush_v net360 net494 VGND VGND VPWR VPWR _01103_ sky130_fd_sc_hd__and3_1
XFILLER_0_88_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_07452_ _01757_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_603 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_07383_ u_decod.rf_ff_res_data_i\[19\] _01550_ _01773_ _02594_ _02614_ VGND VGND
+ VPWR VPWR _02615_ sky130_fd_sc_hd__a221o_1
X_06403_ _01672_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__buf_8
XFILLER_0_134_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_600 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09122_ _04252_ _04254_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__xnor2_1
X_06334_ _01512_ _01515_ _01558_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_33_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_767 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09053_ _04194_ u_exe.branch_v VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__and2_1
X_06265_ u_decod.rf_ff_rd_adr_q_i\[3\] VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_853 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_08004_ _03188_ _03209_ _03198_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__and3_4
X_06196_ _01455_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_897 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_461 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09955_ u_decod.rf_ff_res_data_i\[28\] VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08906_ u_decod.rs1_data_q\[13\] u_decod.branch_imm_q_o\[13\] VGND VGND VPWR VPWR
+ _04068_ sky130_fd_sc_hd__and2_1
X_09886_ _04733_ VGND VGND VPWR VPWR _00229_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_146_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ u_decod.branch_imm_q_o\[0\] _01061_ _01060_ _04002_ _03999_ VGND VGND VPWR
+ VPWR _04009_ sky130_fd_sc_hd__a311o_1
X_08768_ _03937_ _03939_ _03941_ _03943_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__or4_1
XFILLER_0_79_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_07719_ u_rf.reg6_q\[26\] _01557_ _02375_ u_rf.reg11_q\[26\] VGND VGND VPWR VPWR
+ _02937_ sky130_fd_sc_hd__a22o_1
X_08699_ u_rf.reg22_q\[25\] _03409_ _03410_ u_rf.reg3_q\[25\] VGND VGND VPWR VPWR
+ _03878_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_49_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10730_ u_rf.reg18_q\[20\] _04980_ _05210_ VGND VGND VPWR VPWR _05211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10661_ _05151_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__buf_6
XFILLER_0_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12400_ clknet_leaf_36_clk _00437_ net273 VGND VGND VPWR VPWR u_rf.reg13_q\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10592_ _05137_ VGND VGND VPWR VPWR _00531_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_11_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12331_ clknet_leaf_136_clk _00368_ net205 VGND VGND VPWR VPWR u_rf.reg11_q\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_236 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12262_ clknet_leaf_139_clk _00299_ net202 VGND VGND VPWR VPWR u_rf.reg9_q\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_11213_ u_rf.reg25_q\[23\] _04987_ _05463_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_157 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12193_ clknet_leaf_117_clk _00230_ net325 VGND VGND VPWR VPWR u_rf.reg7_q\[6\] sky130_fd_sc_hd__dfrtp_1
X_11144_ _05430_ VGND VGND VPWR VPWR _00790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_11075_ _04768_ u_rf.reg23_q\[22\] _05391_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_393 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10026_ u_rf.reg8_q\[27\] _04484_ _04812_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11977_ clknet_leaf_77_clk net464 net369 VGND VGND VPWR VPWR u_decod.pc_q_o\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_19_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10928_ u_rf.reg21_q\[17\] _04974_ _05308_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_533 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10859_ u_rf.reg20_q\[17\] _04974_ _05271_ VGND VGND VPWR VPWR _05279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12529_ clknet_leaf_55_clk _00566_ net296 VGND VGND VPWR VPWR u_rf.reg17_q\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_06050_ _01312_ _01313_ _01319_ _01320_ VGND VGND VPWR VPWR _01321_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_41_258 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_45 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_645 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout308 net309 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__buf_4
Xfanout319 net320 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_4
X_06952_ _01442_ _02188_ _02195_ _02200_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a31o_1
X_09740_ _04652_ VGND VGND VPWR VPWR _00164_ sky130_fd_sc_hd__clkbuf_1
.ends

